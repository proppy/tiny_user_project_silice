magic
tech sky130A
magscale 1 2
timestamp 1671820187
<< viali >>
rect 6009 31433 6043 31467
rect 13645 31433 13679 31467
rect 2320 31365 2354 31399
rect 9229 31365 9263 31399
rect 14556 31365 14590 31399
rect 19441 31365 19475 31399
rect 19657 31365 19691 31399
rect 4169 31297 4203 31331
rect 4629 31297 4663 31331
rect 4896 31297 4930 31331
rect 6561 31297 6595 31331
rect 6745 31297 6779 31331
rect 7205 31297 7239 31331
rect 7472 31297 7506 31331
rect 9321 31297 9355 31331
rect 10048 31297 10082 31331
rect 12837 31297 12871 31331
rect 14289 31297 14323 31331
rect 16129 31297 16163 31331
rect 17121 31297 17155 31331
rect 18705 31297 18739 31331
rect 20269 31297 20303 31331
rect 20453 31297 20487 31331
rect 20545 31297 20579 31331
rect 21005 31297 21039 31331
rect 22017 31297 22051 31331
rect 23857 31297 23891 31331
rect 24961 31297 24995 31331
rect 27169 31297 27203 31331
rect 28181 31297 28215 31331
rect 2053 31229 2087 31263
rect 9781 31229 9815 31263
rect 13093 31229 13127 31263
rect 16865 31229 16899 31263
rect 3433 31161 3467 31195
rect 11713 31161 11747 31195
rect 18245 31161 18279 31195
rect 19809 31161 19843 31195
rect 4077 31093 4111 31127
rect 6745 31093 6779 31127
rect 8585 31093 8619 31127
rect 11161 31093 11195 31127
rect 15669 31093 15703 31127
rect 19625 31093 19659 31127
rect 20269 31093 20303 31127
rect 8585 30889 8619 30923
rect 18245 30889 18279 30923
rect 21373 30889 21407 30923
rect 27721 30889 27755 30923
rect 28365 30889 28399 30923
rect 4905 30821 4939 30855
rect 11161 30821 11195 30855
rect 11621 30821 11655 30855
rect 18061 30821 18095 30855
rect 19441 30821 19475 30855
rect 12265 30753 12299 30787
rect 15669 30753 15703 30787
rect 19717 30753 19751 30787
rect 20821 30753 20855 30787
rect 2053 30685 2087 30719
rect 4353 30685 4387 30719
rect 6489 30685 6523 30719
rect 6745 30685 6779 30719
rect 7205 30685 7239 30719
rect 9137 30685 9171 30719
rect 9321 30685 9355 30719
rect 9781 30685 9815 30719
rect 12532 30685 12566 30719
rect 15402 30685 15436 30719
rect 17141 30685 17175 30719
rect 17325 30685 17359 30719
rect 17509 30685 17543 30719
rect 17601 30685 17635 30719
rect 19441 30685 19475 30719
rect 19533 30685 19567 30719
rect 20177 30685 20211 30719
rect 20361 30685 20395 30719
rect 2320 30617 2354 30651
rect 4537 30617 4571 30651
rect 4629 30617 4663 30651
rect 7472 30617 7506 30651
rect 10048 30617 10082 30651
rect 16681 30617 16715 30651
rect 18429 30617 18463 30651
rect 3433 30549 3467 30583
rect 4721 30549 4755 30583
rect 5365 30549 5399 30583
rect 9229 30549 9263 30583
rect 13645 30549 13679 30583
rect 14289 30549 14323 30583
rect 16129 30549 16163 30583
rect 16313 30549 16347 30583
rect 16405 30549 16439 30583
rect 16497 30549 16531 30583
rect 18229 30549 18263 30583
rect 20269 30549 20303 30583
rect 10885 30345 10919 30379
rect 15761 30345 15795 30379
rect 19993 30345 20027 30379
rect 3056 30277 3090 30311
rect 6653 30277 6687 30311
rect 14688 30277 14722 30311
rect 15577 30277 15611 30311
rect 15669 30277 15703 30311
rect 19441 30277 19475 30311
rect 20545 30277 20579 30311
rect 2053 30209 2087 30243
rect 2329 30209 2363 30243
rect 4629 30209 4663 30243
rect 4896 30209 4930 30243
rect 6552 30209 6586 30243
rect 6833 30209 6867 30243
rect 7921 30209 7955 30243
rect 9761 30209 9795 30243
rect 11969 30209 12003 30243
rect 14933 30209 14967 30243
rect 15393 30209 15427 30243
rect 17141 30209 17175 30243
rect 17969 30209 18003 30243
rect 18613 30209 18647 30243
rect 19349 30209 19383 30243
rect 19533 30209 19567 30243
rect 2237 30141 2271 30175
rect 2789 30141 2823 30175
rect 7665 30141 7699 30175
rect 9505 30141 9539 30175
rect 11713 30141 11747 30175
rect 16865 30141 16899 30175
rect 18153 30141 18187 30175
rect 1869 30073 1903 30107
rect 4169 30073 4203 30107
rect 6009 30073 6043 30107
rect 18797 30073 18831 30107
rect 6837 30005 6871 30039
rect 9045 30005 9079 30039
rect 13093 30005 13127 30039
rect 13553 30005 13587 30039
rect 15945 30005 15979 30039
rect 16957 30005 16991 30039
rect 17325 30005 17359 30039
rect 17785 30005 17819 30039
rect 28365 30005 28399 30039
rect 15301 29801 15335 29835
rect 17325 29801 17359 29835
rect 4905 29733 4939 29767
rect 7205 29733 7239 29767
rect 11713 29733 11747 29767
rect 13645 29733 13679 29767
rect 15669 29733 15703 29767
rect 18245 29733 18279 29767
rect 18705 29733 18739 29767
rect 13093 29665 13127 29699
rect 14841 29665 14875 29699
rect 2053 29597 2087 29631
rect 4537 29597 4571 29631
rect 6745 29597 6779 29631
rect 8585 29597 8619 29631
rect 9413 29597 9447 29631
rect 14289 29597 14323 29631
rect 14473 29597 14507 29631
rect 14565 29597 14599 29631
rect 15485 29597 15519 29631
rect 15761 29597 15795 29631
rect 16221 29597 16255 29631
rect 16405 29597 16439 29631
rect 16589 29597 16623 29631
rect 16681 29597 16715 29631
rect 17969 29597 18003 29631
rect 18705 29597 18739 29631
rect 18889 29597 18923 29631
rect 28365 29597 28399 29631
rect 2320 29529 2354 29563
rect 4353 29529 4387 29563
rect 4721 29529 4755 29563
rect 6500 29529 6534 29563
rect 8340 29529 8374 29563
rect 9680 29529 9714 29563
rect 12848 29529 12882 29563
rect 17509 29529 17543 29563
rect 18245 29529 18279 29563
rect 19441 29529 19475 29563
rect 19993 29529 20027 29563
rect 20545 29529 20579 29563
rect 3433 29461 3467 29495
rect 4629 29461 4663 29495
rect 5365 29461 5399 29495
rect 10793 29461 10827 29495
rect 14657 29461 14691 29495
rect 17141 29461 17175 29495
rect 17309 29461 17343 29495
rect 18061 29461 18095 29495
rect 2329 29257 2363 29291
rect 6009 29257 6043 29291
rect 8309 29257 8343 29291
rect 11805 29257 11839 29291
rect 12449 29257 12483 29291
rect 16037 29257 16071 29291
rect 17049 29257 17083 29291
rect 1961 29121 1995 29155
rect 2145 29121 2179 29155
rect 2789 29121 2823 29155
rect 3056 29121 3090 29155
rect 4629 29121 4663 29155
rect 4896 29121 4930 29155
rect 6561 29121 6595 29155
rect 9597 29121 9631 29155
rect 10057 29121 10091 29155
rect 12265 29121 12299 29155
rect 13001 29121 13035 29155
rect 14749 29121 14783 29155
rect 15577 29121 15611 29155
rect 15669 29121 15703 29155
rect 15853 29121 15887 29155
rect 16865 29121 16899 29155
rect 17141 29121 17175 29155
rect 17601 29121 17635 29155
rect 17785 29121 17819 29155
rect 18245 29121 18279 29155
rect 1869 29053 1903 29087
rect 6837 29053 6871 29087
rect 4169 28985 4203 29019
rect 11161 28985 11195 29019
rect 16865 28985 16899 29019
rect 17601 28985 17635 29019
rect 5549 28713 5583 28747
rect 8493 28713 8527 28747
rect 11345 28713 11379 28747
rect 14289 28713 14323 28747
rect 15393 28713 15427 28747
rect 15761 28713 15795 28747
rect 16497 28713 16531 28747
rect 3433 28645 3467 28679
rect 8033 28645 8067 28679
rect 9735 28645 9769 28679
rect 17049 28645 17083 28679
rect 18245 28645 18279 28679
rect 7481 28577 7515 28611
rect 9965 28577 9999 28611
rect 13645 28577 13679 28611
rect 14448 28577 14482 28611
rect 14565 28577 14599 28611
rect 14657 28577 14691 28611
rect 14933 28577 14967 28611
rect 15853 28577 15887 28611
rect 16405 28577 16439 28611
rect 16589 28577 16623 28611
rect 2053 28509 2087 28543
rect 4813 28509 4847 28543
rect 7021 28509 7055 28543
rect 13277 28509 13311 28543
rect 13461 28509 13495 28543
rect 15577 28509 15611 28543
rect 16313 28509 16347 28543
rect 17049 28509 17083 28543
rect 17233 28509 17267 28543
rect 17693 28509 17727 28543
rect 2320 28441 2354 28475
rect 4169 28441 4203 28475
rect 7665 28441 7699 28475
rect 12633 28441 12667 28475
rect 7757 28373 7791 28407
rect 7849 28373 7883 28407
rect 13093 28373 13127 28407
rect 13369 28373 13403 28407
rect 8953 28169 8987 28203
rect 10793 28169 10827 28203
rect 3188 28101 3222 28135
rect 9680 28101 9714 28135
rect 14841 28101 14875 28135
rect 3433 28033 3467 28067
rect 4077 28033 4111 28067
rect 4629 28033 4663 28067
rect 4896 28033 4930 28067
rect 6745 28033 6779 28067
rect 7573 28033 7607 28067
rect 7829 28033 7863 28067
rect 9413 28033 9447 28067
rect 11980 28033 12014 28067
rect 14105 28033 14139 28067
rect 15025 28033 15059 28067
rect 15853 28033 15887 28067
rect 15945 28033 15979 28067
rect 6837 27965 6871 27999
rect 6929 27965 6963 27999
rect 7021 27965 7055 27999
rect 11713 27965 11747 27999
rect 14381 27965 14415 27999
rect 15301 27965 15335 27999
rect 3893 27897 3927 27931
rect 6561 27897 6595 27931
rect 16865 27897 16899 27931
rect 2053 27829 2087 27863
rect 6009 27829 6043 27863
rect 13093 27829 13127 27863
rect 13921 27829 13955 27863
rect 14289 27829 14323 27863
rect 15209 27829 15243 27863
rect 16129 27829 16163 27863
rect 28365 27829 28399 27863
rect 4353 27625 4387 27659
rect 15301 27625 15335 27659
rect 3433 27557 3467 27591
rect 5365 27557 5399 27591
rect 11253 27557 11287 27591
rect 15945 27557 15979 27591
rect 16681 27557 16715 27591
rect 1961 27489 1995 27523
rect 4825 27489 4859 27523
rect 10701 27489 10735 27523
rect 12541 27489 12575 27523
rect 13369 27489 13403 27523
rect 2145 27421 2179 27455
rect 3341 27421 3375 27455
rect 3433 27421 3467 27455
rect 4537 27421 4571 27455
rect 4721 27421 4755 27455
rect 6745 27421 6779 27455
rect 7205 27421 7239 27455
rect 10445 27421 10479 27455
rect 12265 27421 12299 27455
rect 13185 27421 13219 27455
rect 13461 27421 13495 27455
rect 16129 27421 16163 27455
rect 16221 27421 16255 27455
rect 16681 27421 16715 27455
rect 16865 27421 16899 27455
rect 28365 27421 28399 27455
rect 3157 27353 3191 27387
rect 6478 27353 6512 27387
rect 7450 27353 7484 27387
rect 14473 27353 14507 27387
rect 14657 27353 14691 27387
rect 15485 27353 15519 27387
rect 15945 27353 15979 27387
rect 17325 27353 17359 27387
rect 2329 27285 2363 27319
rect 8585 27285 8619 27319
rect 9321 27285 9355 27319
rect 13001 27285 13035 27319
rect 14289 27285 14323 27319
rect 15117 27285 15151 27319
rect 15285 27285 15319 27319
rect 1685 27081 1719 27115
rect 3249 27081 3283 27115
rect 3985 27081 4019 27115
rect 10609 27081 10643 27115
rect 13001 27081 13035 27115
rect 14841 27081 14875 27115
rect 15669 27081 15703 27115
rect 16221 27081 16255 27115
rect 5764 27013 5798 27047
rect 8769 27013 8803 27047
rect 11069 27013 11103 27047
rect 13921 27013 13955 27047
rect 14121 27013 14155 27047
rect 1869 26945 1903 26979
rect 2605 26945 2639 26979
rect 3157 26945 3191 26979
rect 3433 26945 3467 26979
rect 3893 26945 3927 26979
rect 4077 26945 4111 26979
rect 6009 26945 6043 26979
rect 7674 26945 7708 26979
rect 7941 26945 7975 26979
rect 8585 26945 8619 26979
rect 9485 26945 9519 26979
rect 13185 26945 13219 26979
rect 13369 26945 13403 26979
rect 14749 26945 14783 26979
rect 15025 26945 15059 26979
rect 15485 26945 15519 26979
rect 8401 26877 8435 26911
rect 9229 26877 9263 26911
rect 12265 26877 12299 26911
rect 12541 26877 12575 26911
rect 13461 26877 13495 26911
rect 2421 26809 2455 26843
rect 14289 26809 14323 26843
rect 15025 26809 15059 26843
rect 3433 26741 3467 26775
rect 4629 26741 4663 26775
rect 6561 26741 6595 26775
rect 14105 26741 14139 26775
rect 2513 26537 2547 26571
rect 4813 26537 4847 26571
rect 5917 26537 5951 26571
rect 7205 26537 7239 26571
rect 12817 26537 12851 26571
rect 13001 26537 13035 26571
rect 3249 26469 3283 26503
rect 4169 26469 4203 26503
rect 5549 26469 5583 26503
rect 6469 26469 6503 26503
rect 8401 26469 8435 26503
rect 13737 26469 13771 26503
rect 6561 26401 6595 26435
rect 8585 26401 8619 26435
rect 9137 26401 9171 26435
rect 11161 26401 11195 26435
rect 11713 26401 11747 26435
rect 12081 26401 12115 26435
rect 13645 26401 13679 26435
rect 1593 26333 1627 26367
rect 2237 26333 2271 26367
rect 3157 26333 3191 26367
rect 3249 26333 3283 26367
rect 3985 26333 4019 26367
rect 4169 26333 4203 26367
rect 4629 26333 4663 26367
rect 5733 26333 5767 26367
rect 6009 26333 6043 26367
rect 6469 26333 6503 26367
rect 7757 26333 7791 26367
rect 8309 26333 8343 26367
rect 11897 26333 11931 26367
rect 12173 26333 12207 26367
rect 13737 26333 13771 26367
rect 14289 26333 14323 26367
rect 14473 26333 14507 26367
rect 2513 26265 2547 26299
rect 2973 26265 3007 26299
rect 6745 26265 6779 26299
rect 8585 26265 8619 26299
rect 9382 26265 9416 26299
rect 12633 26265 12667 26299
rect 12849 26265 12883 26299
rect 13461 26265 13495 26299
rect 14933 26265 14967 26299
rect 2329 26197 2363 26231
rect 10517 26197 10551 26231
rect 14381 26197 14415 26231
rect 15485 26197 15519 26231
rect 1685 25993 1719 26027
rect 7205 25993 7239 26027
rect 8309 25993 8343 26027
rect 10517 25993 10551 26027
rect 10977 25993 11011 26027
rect 12801 25993 12835 26027
rect 6009 25925 6043 25959
rect 6561 25925 6595 25959
rect 9597 25925 9631 25959
rect 11713 25925 11747 25959
rect 13001 25925 13035 25959
rect 14749 25925 14783 25959
rect 1869 25857 1903 25891
rect 3985 25857 4019 25891
rect 5733 25857 5767 25891
rect 5825 25857 5859 25891
rect 7113 25857 7147 25891
rect 7389 25857 7423 25891
rect 10057 25857 10091 25891
rect 10333 25857 10367 25891
rect 11897 25857 11931 25891
rect 13449 25857 13483 25891
rect 13645 25857 13679 25891
rect 17141 25857 17175 25891
rect 17601 25857 17635 25891
rect 2973 25789 3007 25823
rect 5089 25789 5123 25823
rect 12173 25789 12207 25823
rect 14105 25789 14139 25823
rect 6009 25721 6043 25755
rect 7389 25721 7423 25755
rect 16957 25721 16991 25755
rect 28365 25721 28399 25755
rect 2329 25653 2363 25687
rect 10149 25653 10183 25687
rect 12081 25653 12115 25687
rect 12633 25653 12667 25687
rect 12817 25653 12851 25687
rect 13645 25653 13679 25687
rect 2237 25449 2271 25483
rect 7389 25449 7423 25483
rect 8217 25449 8251 25483
rect 8585 25449 8619 25483
rect 10149 25449 10183 25483
rect 12725 25449 12759 25483
rect 1593 25381 1627 25415
rect 4905 25381 4939 25415
rect 6009 25381 6043 25415
rect 6929 25381 6963 25415
rect 28365 25381 28399 25415
rect 6837 25313 6871 25347
rect 8125 25313 8159 25347
rect 6193 25245 6227 25279
rect 6929 25245 6963 25279
rect 7665 25245 7699 25279
rect 8401 25245 8435 25279
rect 9873 25245 9907 25279
rect 9965 25245 9999 25279
rect 10793 25245 10827 25279
rect 10977 25245 11011 25279
rect 11713 25245 11747 25279
rect 11897 25245 11931 25279
rect 13277 25245 13311 25279
rect 3433 25177 3467 25211
rect 5549 25177 5583 25211
rect 6653 25177 6687 25211
rect 7389 25177 7423 25211
rect 12633 25177 12667 25211
rect 4261 25109 4295 25143
rect 7573 25109 7607 25143
rect 9137 25109 9171 25143
rect 10609 25109 10643 25143
rect 12081 25109 12115 25143
rect 14289 25109 14323 25143
rect 2145 24905 2179 24939
rect 8217 24837 8251 24871
rect 9597 24837 9631 24871
rect 9367 24803 9401 24837
rect 3341 24769 3375 24803
rect 5181 24769 5215 24803
rect 6745 24769 6779 24803
rect 6929 24769 6963 24803
rect 7481 24769 7515 24803
rect 8401 24769 8435 24803
rect 8493 24769 8527 24803
rect 10609 24769 10643 24803
rect 11713 24769 11747 24803
rect 11897 24769 11931 24803
rect 11989 24769 12023 24803
rect 12541 24769 12575 24803
rect 13369 24769 13403 24803
rect 2697 24701 2731 24735
rect 3893 24701 3927 24735
rect 4537 24701 4571 24735
rect 6009 24701 6043 24735
rect 10885 24701 10919 24735
rect 6745 24633 6779 24667
rect 7665 24633 7699 24667
rect 10057 24633 10091 24667
rect 10701 24633 10735 24667
rect 11713 24633 11747 24667
rect 9229 24565 9263 24599
rect 9413 24565 9447 24599
rect 10793 24565 10827 24599
rect 2513 24361 2547 24395
rect 4353 24361 4387 24395
rect 8401 24361 8435 24395
rect 9965 24361 9999 24395
rect 10793 24361 10827 24395
rect 12173 24361 12207 24395
rect 9137 24293 9171 24327
rect 10057 24293 10091 24327
rect 7021 24225 7055 24259
rect 10149 24225 10183 24259
rect 1593 24157 1627 24191
rect 8401 24157 8435 24191
rect 8585 24157 8619 24191
rect 9321 24157 9355 24191
rect 9413 24157 9447 24191
rect 9873 24157 9907 24191
rect 10609 24157 10643 24191
rect 10793 24157 10827 24191
rect 28365 24157 28399 24191
rect 5089 24089 5123 24123
rect 9137 24089 9171 24123
rect 11253 24089 11287 24123
rect 6469 24021 6503 24055
rect 7757 24021 7791 24055
rect 4353 23817 4387 23851
rect 6929 23817 6963 23851
rect 9873 23817 9907 23851
rect 10517 23817 10551 23851
rect 9781 23681 9815 23715
rect 9965 23681 9999 23715
rect 8677 23613 8711 23647
rect 9321 23613 9355 23647
rect 10977 23613 11011 23647
rect 1593 23477 1627 23511
rect 9505 23273 9539 23307
rect 28365 23069 28399 23103
rect 1593 22389 1627 22423
rect 28365 21981 28399 22015
rect 1593 21437 1627 21471
rect 28365 21301 28399 21335
rect 1593 20213 1627 20247
rect 28365 19941 28399 19975
rect 1593 19805 1627 19839
rect 28365 19125 28399 19159
rect 1593 18037 1627 18071
rect 1593 17629 1627 17663
rect 28365 17629 28399 17663
rect 28365 16949 28399 16983
rect 1593 15997 1627 16031
rect 28365 15861 28399 15895
rect 1593 15453 1627 15487
rect 28365 14841 28399 14875
rect 1593 14365 1627 14399
rect 28365 13685 28399 13719
rect 1593 13277 1627 13311
rect 28365 13277 28399 13311
rect 1593 12189 1627 12223
rect 1593 11509 1627 11543
rect 28365 11509 28399 11543
rect 28365 11101 28399 11135
rect 1593 10013 1627 10047
rect 28365 9401 28399 9435
rect 1593 9333 1627 9367
rect 28365 9061 28399 9095
rect 1593 7837 1627 7871
rect 28365 7837 28399 7871
rect 1593 7157 1627 7191
rect 28365 6749 28399 6783
rect 1593 6069 1627 6103
rect 28365 5661 28399 5695
rect 1593 5117 1627 5151
rect 28365 4981 28399 5015
rect 28365 4437 28399 4471
rect 28089 4029 28123 4063
rect 28365 4029 28399 4063
rect 1593 3893 1627 3927
rect 28365 3621 28399 3655
rect 1593 3485 1627 3519
rect 28365 2805 28399 2839
<< metal1 >>
rect 12526 31900 12532 31952
rect 12584 31940 12590 31952
rect 14918 31940 14924 31952
rect 12584 31912 14924 31940
rect 12584 31900 12590 31912
rect 14918 31900 14924 31912
rect 14976 31900 14982 31952
rect 13814 31832 13820 31884
rect 13872 31872 13878 31884
rect 16114 31872 16120 31884
rect 13872 31844 16120 31872
rect 13872 31832 13878 31844
rect 16114 31832 16120 31844
rect 16172 31832 16178 31884
rect 12986 31764 12992 31816
rect 13044 31804 13050 31816
rect 16390 31804 16396 31816
rect 13044 31776 16396 31804
rect 13044 31764 13050 31776
rect 16390 31764 16396 31776
rect 16448 31764 16454 31816
rect 9306 31696 9312 31748
rect 9364 31736 9370 31748
rect 13630 31736 13636 31748
rect 9364 31708 13636 31736
rect 9364 31696 9370 31708
rect 13630 31696 13636 31708
rect 13688 31696 13694 31748
rect 14274 31696 14280 31748
rect 14332 31736 14338 31748
rect 19702 31736 19708 31748
rect 14332 31708 19708 31736
rect 14332 31696 14338 31708
rect 19702 31696 19708 31708
rect 19760 31696 19766 31748
rect 4154 31628 4160 31680
rect 4212 31668 4218 31680
rect 6546 31668 6552 31680
rect 4212 31640 6552 31668
rect 4212 31628 4218 31640
rect 6546 31628 6552 31640
rect 6604 31668 6610 31680
rect 7098 31668 7104 31680
rect 6604 31640 7104 31668
rect 6604 31628 6610 31640
rect 7098 31628 7104 31640
rect 7156 31628 7162 31680
rect 8570 31628 8576 31680
rect 8628 31668 8634 31680
rect 14550 31668 14556 31680
rect 8628 31640 14556 31668
rect 8628 31628 8634 31640
rect 14550 31628 14556 31640
rect 14608 31628 14614 31680
rect 1104 31578 29048 31600
rect 1104 31526 7896 31578
rect 7948 31526 7960 31578
rect 8012 31526 8024 31578
rect 8076 31526 8088 31578
rect 8140 31526 8152 31578
rect 8204 31526 14842 31578
rect 14894 31526 14906 31578
rect 14958 31526 14970 31578
rect 15022 31526 15034 31578
rect 15086 31526 15098 31578
rect 15150 31526 21788 31578
rect 21840 31526 21852 31578
rect 21904 31526 21916 31578
rect 21968 31526 21980 31578
rect 22032 31526 22044 31578
rect 22096 31526 28734 31578
rect 28786 31526 28798 31578
rect 28850 31526 28862 31578
rect 28914 31526 28926 31578
rect 28978 31526 28990 31578
rect 29042 31526 29048 31578
rect 1104 31504 29048 31526
rect 5350 31464 5356 31476
rect 2746 31436 5356 31464
rect 2308 31399 2366 31405
rect 2308 31365 2320 31399
rect 2354 31396 2366 31399
rect 2746 31396 2774 31436
rect 5350 31424 5356 31436
rect 5408 31424 5414 31476
rect 5997 31467 6055 31473
rect 5997 31433 6009 31467
rect 6043 31464 6055 31467
rect 11330 31464 11336 31476
rect 6043 31436 11336 31464
rect 6043 31433 6055 31436
rect 5997 31427 6055 31433
rect 11330 31424 11336 31436
rect 11388 31424 11394 31476
rect 13630 31464 13636 31476
rect 13543 31436 13636 31464
rect 13630 31424 13636 31436
rect 13688 31464 13694 31476
rect 14090 31464 14096 31476
rect 13688 31436 14096 31464
rect 13688 31424 13694 31436
rect 14090 31424 14096 31436
rect 14148 31464 14154 31476
rect 14148 31436 19564 31464
rect 14148 31424 14154 31436
rect 5534 31396 5540 31408
rect 2354 31368 2774 31396
rect 4632 31368 5540 31396
rect 2354 31365 2366 31368
rect 2308 31359 2366 31365
rect 4154 31328 4160 31340
rect 4115 31300 4160 31328
rect 4154 31288 4160 31300
rect 4212 31288 4218 31340
rect 4632 31337 4660 31368
rect 5534 31356 5540 31368
rect 5592 31396 5598 31408
rect 9217 31399 9275 31405
rect 5592 31368 7236 31396
rect 5592 31356 5598 31368
rect 4617 31331 4675 31337
rect 4617 31297 4629 31331
rect 4663 31297 4675 31331
rect 4617 31291 4675 31297
rect 4884 31331 4942 31337
rect 4884 31297 4896 31331
rect 4930 31328 4942 31331
rect 5442 31328 5448 31340
rect 4930 31300 5448 31328
rect 4930 31297 4942 31300
rect 4884 31291 4942 31297
rect 5442 31288 5448 31300
rect 5500 31288 5506 31340
rect 6546 31328 6552 31340
rect 6507 31300 6552 31328
rect 6546 31288 6552 31300
rect 6604 31288 6610 31340
rect 7208 31337 7236 31368
rect 9217 31365 9229 31399
rect 9263 31396 9275 31399
rect 14182 31396 14188 31408
rect 9263 31368 14188 31396
rect 9263 31365 9275 31368
rect 9217 31359 9275 31365
rect 14182 31356 14188 31368
rect 14240 31356 14246 31408
rect 14550 31405 14556 31408
rect 14544 31396 14556 31405
rect 14511 31368 14556 31396
rect 14544 31359 14556 31368
rect 14550 31356 14556 31359
rect 14608 31356 14614 31408
rect 17218 31356 17224 31408
rect 17276 31396 17282 31408
rect 19429 31399 19487 31405
rect 17276 31368 18736 31396
rect 17276 31356 17282 31368
rect 6733 31331 6791 31337
rect 6733 31297 6745 31331
rect 6779 31297 6791 31331
rect 6733 31291 6791 31297
rect 7193 31331 7251 31337
rect 7193 31297 7205 31331
rect 7239 31297 7251 31331
rect 7193 31291 7251 31297
rect 7460 31331 7518 31337
rect 7460 31297 7472 31331
rect 7506 31328 7518 31331
rect 9309 31331 9367 31337
rect 7506 31300 9260 31328
rect 7506 31297 7518 31300
rect 7460 31291 7518 31297
rect 2038 31260 2044 31272
rect 1999 31232 2044 31260
rect 2038 31220 2044 31232
rect 2096 31220 2102 31272
rect 6270 31220 6276 31272
rect 6328 31260 6334 31272
rect 6748 31260 6776 31291
rect 6328 31232 6776 31260
rect 9232 31260 9260 31300
rect 9309 31297 9321 31331
rect 9355 31328 9367 31331
rect 9674 31328 9680 31340
rect 9355 31300 9680 31328
rect 9355 31297 9367 31300
rect 9309 31291 9367 31297
rect 9674 31288 9680 31300
rect 9732 31288 9738 31340
rect 10042 31337 10048 31340
rect 10036 31291 10048 31337
rect 10100 31328 10106 31340
rect 12825 31331 12883 31337
rect 10100 31300 10136 31328
rect 10042 31288 10048 31291
rect 10100 31288 10106 31300
rect 12825 31297 12837 31331
rect 12871 31328 12883 31331
rect 12986 31328 12992 31340
rect 12871 31300 12992 31328
rect 12871 31297 12883 31300
rect 12825 31291 12883 31297
rect 12986 31288 12992 31300
rect 13044 31288 13050 31340
rect 14277 31331 14335 31337
rect 14277 31328 14289 31331
rect 13096 31300 14289 31328
rect 13096 31272 13124 31300
rect 14277 31297 14289 31300
rect 14323 31328 14335 31331
rect 15654 31328 15660 31340
rect 14323 31300 15660 31328
rect 14323 31297 14335 31300
rect 14277 31291 14335 31297
rect 15654 31288 15660 31300
rect 15712 31288 15718 31340
rect 16114 31328 16120 31340
rect 16075 31300 16120 31328
rect 16114 31288 16120 31300
rect 16172 31288 16178 31340
rect 16574 31288 16580 31340
rect 16632 31328 16638 31340
rect 18708 31337 18736 31368
rect 19429 31365 19441 31399
rect 19475 31365 19487 31399
rect 19536 31396 19564 31436
rect 19645 31399 19703 31405
rect 19645 31396 19657 31399
rect 19536 31368 19657 31396
rect 19429 31359 19487 31365
rect 19645 31365 19657 31368
rect 19691 31396 19703 31399
rect 21358 31396 21364 31408
rect 19691 31368 21364 31396
rect 19691 31365 19703 31368
rect 19645 31359 19703 31365
rect 17109 31331 17167 31337
rect 17109 31328 17121 31331
rect 16632 31300 17121 31328
rect 16632 31288 16638 31300
rect 17109 31297 17121 31300
rect 17155 31297 17167 31331
rect 17109 31291 17167 31297
rect 18693 31331 18751 31337
rect 18693 31297 18705 31331
rect 18739 31297 18751 31331
rect 18693 31291 18751 31297
rect 9398 31260 9404 31272
rect 9232 31232 9404 31260
rect 6328 31220 6334 31232
rect 9398 31220 9404 31232
rect 9456 31220 9462 31272
rect 9766 31260 9772 31272
rect 9727 31232 9772 31260
rect 9766 31220 9772 31232
rect 9824 31220 9830 31272
rect 11974 31260 11980 31272
rect 10796 31232 11980 31260
rect 3421 31195 3479 31201
rect 3421 31161 3433 31195
rect 3467 31192 3479 31195
rect 3467 31164 4660 31192
rect 3467 31161 3479 31164
rect 3421 31155 3479 31161
rect 3050 31084 3056 31136
rect 3108 31124 3114 31136
rect 3970 31124 3976 31136
rect 3108 31096 3976 31124
rect 3108 31084 3114 31096
rect 3970 31084 3976 31096
rect 4028 31124 4034 31136
rect 4065 31127 4123 31133
rect 4065 31124 4077 31127
rect 4028 31096 4077 31124
rect 4028 31084 4034 31096
rect 4065 31093 4077 31096
rect 4111 31093 4123 31127
rect 4632 31124 4660 31164
rect 6564 31164 7236 31192
rect 6564 31124 6592 31164
rect 6730 31124 6736 31136
rect 4632 31096 6592 31124
rect 6691 31096 6736 31124
rect 4065 31087 4123 31093
rect 6730 31084 6736 31096
rect 6788 31084 6794 31136
rect 7208 31124 7236 31164
rect 8386 31124 8392 31136
rect 7208 31096 8392 31124
rect 8386 31084 8392 31096
rect 8444 31084 8450 31136
rect 8573 31127 8631 31133
rect 8573 31093 8585 31127
rect 8619 31124 8631 31127
rect 10042 31124 10048 31136
rect 8619 31096 10048 31124
rect 8619 31093 8631 31096
rect 8573 31087 8631 31093
rect 10042 31084 10048 31096
rect 10100 31124 10106 31136
rect 10796 31124 10824 31232
rect 11974 31220 11980 31232
rect 12032 31220 12038 31272
rect 13078 31260 13084 31272
rect 13039 31232 13084 31260
rect 13078 31220 13084 31232
rect 13136 31220 13142 31272
rect 15672 31260 15700 31288
rect 16853 31263 16911 31269
rect 16853 31260 16865 31263
rect 15672 31232 16865 31260
rect 16853 31229 16865 31232
rect 16899 31229 16911 31263
rect 16853 31223 16911 31229
rect 17862 31220 17868 31272
rect 17920 31260 17926 31272
rect 19444 31260 19472 31359
rect 21358 31356 21364 31368
rect 21416 31356 21422 31408
rect 20257 31331 20315 31337
rect 20257 31297 20269 31331
rect 20303 31297 20315 31331
rect 20438 31328 20444 31340
rect 20399 31300 20444 31328
rect 20257 31291 20315 31297
rect 17920 31232 19472 31260
rect 17920 31220 17926 31232
rect 19702 31220 19708 31272
rect 19760 31260 19766 31272
rect 20272 31260 20300 31291
rect 20438 31288 20444 31300
rect 20496 31288 20502 31340
rect 20530 31288 20536 31340
rect 20588 31328 20594 31340
rect 20588 31300 20633 31328
rect 20588 31288 20594 31300
rect 20714 31288 20720 31340
rect 20772 31328 20778 31340
rect 20993 31331 21051 31337
rect 20993 31328 21005 31331
rect 20772 31300 21005 31328
rect 20772 31288 20778 31300
rect 20993 31297 21005 31300
rect 21039 31297 21051 31331
rect 20993 31291 21051 31297
rect 21542 31288 21548 31340
rect 21600 31328 21606 31340
rect 22005 31331 22063 31337
rect 22005 31328 22017 31331
rect 21600 31300 22017 31328
rect 21600 31288 21606 31300
rect 22005 31297 22017 31300
rect 22051 31297 22063 31331
rect 22005 31291 22063 31297
rect 23750 31288 23756 31340
rect 23808 31328 23814 31340
rect 23845 31331 23903 31337
rect 23845 31328 23857 31331
rect 23808 31300 23857 31328
rect 23808 31288 23814 31300
rect 23845 31297 23857 31300
rect 23891 31297 23903 31331
rect 23845 31291 23903 31297
rect 24854 31288 24860 31340
rect 24912 31328 24918 31340
rect 24949 31331 25007 31337
rect 24949 31328 24961 31331
rect 24912 31300 24961 31328
rect 24912 31288 24918 31300
rect 24949 31297 24961 31300
rect 24995 31297 25007 31331
rect 24949 31291 25007 31297
rect 27062 31288 27068 31340
rect 27120 31328 27126 31340
rect 27157 31331 27215 31337
rect 27157 31328 27169 31331
rect 27120 31300 27169 31328
rect 27120 31288 27126 31300
rect 27157 31297 27169 31300
rect 27203 31297 27215 31331
rect 28166 31328 28172 31340
rect 28127 31300 28172 31328
rect 27157 31291 27215 31297
rect 28166 31288 28172 31300
rect 28224 31288 28230 31340
rect 19760 31232 20300 31260
rect 19760 31220 19766 31232
rect 11701 31195 11759 31201
rect 11701 31161 11713 31195
rect 11747 31192 11759 31195
rect 12066 31192 12072 31204
rect 11747 31164 12072 31192
rect 11747 31161 11759 31164
rect 11701 31155 11759 31161
rect 12066 31152 12072 31164
rect 12124 31152 12130 31204
rect 17954 31152 17960 31204
rect 18012 31192 18018 31204
rect 18233 31195 18291 31201
rect 18233 31192 18245 31195
rect 18012 31164 18245 31192
rect 18012 31152 18018 31164
rect 18233 31161 18245 31164
rect 18279 31161 18291 31195
rect 19797 31195 19855 31201
rect 19797 31192 19809 31195
rect 18233 31155 18291 31161
rect 19444 31164 19809 31192
rect 10100 31096 10824 31124
rect 10100 31084 10106 31096
rect 11054 31084 11060 31136
rect 11112 31124 11118 31136
rect 11149 31127 11207 31133
rect 11149 31124 11161 31127
rect 11112 31096 11161 31124
rect 11112 31084 11118 31096
rect 11149 31093 11161 31096
rect 11195 31093 11207 31127
rect 11149 31087 11207 31093
rect 11330 31084 11336 31136
rect 11388 31124 11394 31136
rect 13446 31124 13452 31136
rect 11388 31096 13452 31124
rect 11388 31084 11394 31096
rect 13446 31084 13452 31096
rect 13504 31084 13510 31136
rect 13906 31084 13912 31136
rect 13964 31124 13970 31136
rect 15562 31124 15568 31136
rect 13964 31096 15568 31124
rect 13964 31084 13970 31096
rect 15562 31084 15568 31096
rect 15620 31084 15626 31136
rect 15657 31127 15715 31133
rect 15657 31093 15669 31127
rect 15703 31124 15715 31127
rect 18046 31124 18052 31136
rect 15703 31096 18052 31124
rect 15703 31093 15715 31096
rect 15657 31087 15715 31093
rect 18046 31084 18052 31096
rect 18104 31084 18110 31136
rect 18138 31084 18144 31136
rect 18196 31124 18202 31136
rect 19444 31124 19472 31164
rect 19797 31161 19809 31164
rect 19843 31192 19855 31195
rect 20162 31192 20168 31204
rect 19843 31164 20168 31192
rect 19843 31161 19855 31164
rect 19797 31155 19855 31161
rect 20162 31152 20168 31164
rect 20220 31152 20226 31204
rect 19610 31124 19616 31136
rect 18196 31096 19472 31124
rect 19571 31096 19616 31124
rect 18196 31084 18202 31096
rect 19610 31084 19616 31096
rect 19668 31084 19674 31136
rect 19886 31084 19892 31136
rect 19944 31124 19950 31136
rect 20257 31127 20315 31133
rect 20257 31124 20269 31127
rect 19944 31096 20269 31124
rect 19944 31084 19950 31096
rect 20257 31093 20269 31096
rect 20303 31093 20315 31127
rect 20257 31087 20315 31093
rect 1104 31034 28888 31056
rect 1104 30982 4423 31034
rect 4475 30982 4487 31034
rect 4539 30982 4551 31034
rect 4603 30982 4615 31034
rect 4667 30982 4679 31034
rect 4731 30982 11369 31034
rect 11421 30982 11433 31034
rect 11485 30982 11497 31034
rect 11549 30982 11561 31034
rect 11613 30982 11625 31034
rect 11677 30982 18315 31034
rect 18367 30982 18379 31034
rect 18431 30982 18443 31034
rect 18495 30982 18507 31034
rect 18559 30982 18571 31034
rect 18623 30982 25261 31034
rect 25313 30982 25325 31034
rect 25377 30982 25389 31034
rect 25441 30982 25453 31034
rect 25505 30982 25517 31034
rect 25569 30982 28888 31034
rect 1104 30960 28888 30982
rect 7190 30920 7196 30932
rect 4908 30892 7196 30920
rect 4908 30861 4936 30892
rect 7190 30880 7196 30892
rect 7248 30880 7254 30932
rect 8570 30920 8576 30932
rect 8531 30892 8576 30920
rect 8570 30880 8576 30892
rect 8628 30880 8634 30932
rect 9766 30880 9772 30932
rect 9824 30920 9830 30932
rect 12986 30920 12992 30932
rect 9824 30892 12992 30920
rect 9824 30880 9830 30892
rect 4893 30855 4951 30861
rect 4893 30821 4905 30855
rect 4939 30821 4951 30855
rect 4893 30815 4951 30821
rect 11149 30855 11207 30861
rect 11149 30821 11161 30855
rect 11195 30821 11207 30855
rect 11149 30815 11207 30821
rect 4706 30744 4712 30796
rect 4764 30784 4770 30796
rect 5074 30784 5080 30796
rect 4764 30756 5080 30784
rect 4764 30744 4770 30756
rect 5074 30744 5080 30756
rect 5132 30744 5138 30796
rect 11164 30784 11192 30815
rect 11330 30812 11336 30864
rect 11388 30852 11394 30864
rect 11609 30855 11667 30861
rect 11609 30852 11621 30855
rect 11388 30824 11621 30852
rect 11388 30812 11394 30824
rect 11609 30821 11621 30824
rect 11655 30821 11667 30855
rect 11609 30815 11667 30821
rect 12158 30784 12164 30796
rect 11164 30756 12164 30784
rect 12158 30744 12164 30756
rect 12216 30744 12222 30796
rect 12268 30793 12296 30892
rect 12986 30880 12992 30892
rect 13044 30880 13050 30932
rect 14182 30880 14188 30932
rect 14240 30920 14246 30932
rect 18233 30923 18291 30929
rect 18233 30920 18245 30923
rect 14240 30892 18245 30920
rect 14240 30880 14246 30892
rect 18233 30889 18245 30892
rect 18279 30920 18291 30923
rect 20438 30920 20444 30932
rect 18279 30892 20444 30920
rect 18279 30889 18291 30892
rect 18233 30883 18291 30889
rect 20438 30880 20444 30892
rect 20496 30880 20502 30932
rect 21358 30920 21364 30932
rect 21319 30892 21364 30920
rect 21358 30880 21364 30892
rect 21416 30880 21422 30932
rect 27706 30920 27712 30932
rect 27667 30892 27712 30920
rect 27706 30880 27712 30892
rect 27764 30880 27770 30932
rect 28350 30920 28356 30932
rect 28311 30892 28356 30920
rect 28350 30880 28356 30892
rect 28408 30880 28414 30932
rect 13354 30812 13360 30864
rect 13412 30852 13418 30864
rect 14550 30852 14556 30864
rect 13412 30824 14556 30852
rect 13412 30812 13418 30824
rect 14550 30812 14556 30824
rect 14608 30812 14614 30864
rect 16114 30812 16120 30864
rect 16172 30852 16178 30864
rect 18049 30855 18107 30861
rect 18049 30852 18061 30855
rect 16172 30824 18061 30852
rect 16172 30812 16178 30824
rect 18049 30821 18061 30824
rect 18095 30821 18107 30855
rect 18049 30815 18107 30821
rect 18782 30812 18788 30864
rect 18840 30852 18846 30864
rect 19429 30855 19487 30861
rect 18840 30824 19380 30852
rect 18840 30812 18846 30824
rect 12253 30787 12311 30793
rect 12253 30753 12265 30787
rect 12299 30753 12311 30787
rect 12253 30747 12311 30753
rect 13262 30744 13268 30796
rect 13320 30784 13326 30796
rect 13998 30784 14004 30796
rect 13320 30756 14004 30784
rect 13320 30744 13326 30756
rect 13998 30744 14004 30756
rect 14056 30744 14062 30796
rect 15654 30784 15660 30796
rect 15615 30756 15660 30784
rect 15654 30744 15660 30756
rect 15712 30744 15718 30796
rect 16850 30744 16856 30796
rect 16908 30784 16914 30796
rect 19242 30784 19248 30796
rect 16908 30756 19248 30784
rect 16908 30744 16914 30756
rect 19242 30744 19248 30756
rect 19300 30744 19306 30796
rect 19352 30784 19380 30824
rect 19429 30821 19441 30855
rect 19475 30852 19487 30855
rect 19794 30852 19800 30864
rect 19475 30824 19800 30852
rect 19475 30821 19487 30824
rect 19429 30815 19487 30821
rect 19794 30812 19800 30824
rect 19852 30812 19858 30864
rect 19705 30787 19763 30793
rect 19705 30784 19717 30787
rect 19352 30756 19717 30784
rect 19705 30753 19717 30756
rect 19751 30784 19763 30787
rect 20809 30787 20867 30793
rect 20809 30784 20821 30787
rect 19751 30756 20821 30784
rect 19751 30753 19763 30756
rect 19705 30747 19763 30753
rect 20809 30753 20821 30756
rect 20855 30753 20867 30787
rect 20809 30747 20867 30753
rect 2038 30716 2044 30728
rect 1951 30688 2044 30716
rect 2038 30676 2044 30688
rect 2096 30716 2102 30728
rect 2682 30716 2688 30728
rect 2096 30688 2688 30716
rect 2096 30676 2102 30688
rect 2682 30676 2688 30688
rect 2740 30676 2746 30728
rect 4341 30719 4399 30725
rect 4341 30685 4353 30719
rect 4387 30716 4399 30719
rect 6178 30716 6184 30728
rect 4387 30688 6184 30716
rect 4387 30685 4399 30688
rect 4341 30679 4399 30685
rect 6178 30676 6184 30688
rect 6236 30676 6242 30728
rect 6477 30719 6535 30725
rect 6477 30685 6489 30719
rect 6523 30716 6535 30719
rect 6638 30716 6644 30728
rect 6523 30688 6644 30716
rect 6523 30685 6535 30688
rect 6477 30679 6535 30685
rect 6638 30676 6644 30688
rect 6696 30676 6702 30728
rect 6733 30719 6791 30725
rect 6733 30685 6745 30719
rect 6779 30716 6791 30719
rect 7193 30719 7251 30725
rect 7193 30716 7205 30719
rect 6779 30688 7205 30716
rect 6779 30685 6791 30688
rect 6733 30679 6791 30685
rect 7193 30685 7205 30688
rect 7239 30716 7251 30719
rect 9125 30719 9183 30725
rect 7239 30688 7696 30716
rect 7239 30685 7251 30688
rect 7193 30679 7251 30685
rect 7668 30660 7696 30688
rect 9125 30685 9137 30719
rect 9171 30716 9183 30719
rect 9214 30716 9220 30728
rect 9171 30688 9220 30716
rect 9171 30685 9183 30688
rect 9125 30679 9183 30685
rect 9214 30676 9220 30688
rect 9272 30676 9278 30728
rect 9306 30676 9312 30728
rect 9364 30716 9370 30728
rect 9769 30719 9827 30725
rect 9364 30688 9457 30716
rect 9364 30676 9370 30688
rect 9769 30685 9781 30719
rect 9815 30716 9827 30719
rect 10962 30716 10968 30728
rect 9815 30688 10968 30716
rect 9815 30685 9827 30688
rect 9769 30679 9827 30685
rect 10962 30676 10968 30688
rect 11020 30676 11026 30728
rect 12520 30719 12578 30725
rect 11072 30688 12434 30716
rect 2308 30651 2366 30657
rect 2308 30617 2320 30651
rect 2354 30648 2366 30651
rect 4062 30648 4068 30660
rect 2354 30620 4068 30648
rect 2354 30617 2366 30620
rect 2308 30611 2366 30617
rect 4062 30608 4068 30620
rect 4120 30608 4126 30660
rect 4246 30608 4252 30660
rect 4304 30648 4310 30660
rect 4525 30651 4583 30657
rect 4525 30648 4537 30651
rect 4304 30620 4537 30648
rect 4304 30608 4310 30620
rect 4525 30617 4537 30620
rect 4571 30617 4583 30651
rect 4525 30611 4583 30617
rect 4617 30651 4675 30657
rect 4617 30617 4629 30651
rect 4663 30648 4675 30651
rect 7460 30651 7518 30657
rect 4663 30620 7420 30648
rect 4663 30617 4675 30620
rect 4617 30611 4675 30617
rect 3421 30583 3479 30589
rect 3421 30549 3433 30583
rect 3467 30580 3479 30583
rect 4338 30580 4344 30592
rect 3467 30552 4344 30580
rect 3467 30549 3479 30552
rect 3421 30543 3479 30549
rect 4338 30540 4344 30552
rect 4396 30540 4402 30592
rect 4706 30580 4712 30592
rect 4667 30552 4712 30580
rect 4706 30540 4712 30552
rect 4764 30540 4770 30592
rect 5353 30583 5411 30589
rect 5353 30549 5365 30583
rect 5399 30580 5411 30583
rect 7282 30580 7288 30592
rect 5399 30552 7288 30580
rect 5399 30549 5411 30552
rect 5353 30543 5411 30549
rect 7282 30540 7288 30552
rect 7340 30540 7346 30592
rect 7392 30580 7420 30620
rect 7460 30617 7472 30651
rect 7506 30648 7518 30651
rect 7558 30648 7564 30660
rect 7506 30620 7564 30648
rect 7506 30617 7518 30620
rect 7460 30611 7518 30617
rect 7558 30608 7564 30620
rect 7616 30608 7622 30660
rect 7650 30608 7656 30660
rect 7708 30608 7714 30660
rect 9324 30648 9352 30676
rect 9140 30620 9352 30648
rect 10036 30651 10094 30657
rect 9140 30580 9168 30620
rect 10036 30617 10048 30651
rect 10082 30648 10094 30651
rect 10594 30648 10600 30660
rect 10082 30620 10600 30648
rect 10082 30617 10094 30620
rect 10036 30611 10094 30617
rect 10594 30608 10600 30620
rect 10652 30608 10658 30660
rect 11072 30648 11100 30688
rect 10796 30620 11100 30648
rect 12406 30648 12434 30688
rect 12520 30685 12532 30719
rect 12566 30716 12578 30719
rect 15102 30716 15108 30728
rect 12566 30688 15108 30716
rect 12566 30685 12578 30688
rect 12520 30679 12578 30685
rect 15102 30676 15108 30688
rect 15160 30676 15166 30728
rect 15378 30676 15384 30728
rect 15436 30725 15442 30728
rect 15436 30716 15448 30725
rect 17129 30719 17187 30725
rect 17129 30716 17141 30719
rect 15436 30688 15481 30716
rect 15548 30688 17141 30716
rect 15436 30679 15448 30688
rect 15436 30676 15442 30679
rect 13262 30648 13268 30660
rect 12406 30620 13268 30648
rect 7392 30552 9168 30580
rect 9217 30583 9275 30589
rect 9217 30549 9229 30583
rect 9263 30580 9275 30583
rect 10796 30580 10824 30620
rect 13262 30608 13268 30620
rect 13320 30608 13326 30660
rect 13372 30620 14320 30648
rect 9263 30552 10824 30580
rect 9263 30549 9275 30552
rect 9217 30543 9275 30549
rect 10870 30540 10876 30592
rect 10928 30580 10934 30592
rect 13372 30580 13400 30620
rect 13630 30580 13636 30592
rect 10928 30552 13400 30580
rect 13591 30552 13636 30580
rect 10928 30540 10934 30552
rect 13630 30540 13636 30552
rect 13688 30540 13694 30592
rect 14292 30589 14320 30620
rect 14550 30608 14556 30660
rect 14608 30648 14614 30660
rect 15548 30648 15576 30688
rect 17129 30685 17141 30688
rect 17175 30685 17187 30719
rect 17310 30716 17316 30728
rect 17271 30688 17316 30716
rect 17129 30679 17187 30685
rect 17310 30676 17316 30688
rect 17368 30676 17374 30728
rect 17494 30716 17500 30728
rect 17455 30688 17500 30716
rect 17494 30676 17500 30688
rect 17552 30676 17558 30728
rect 17604 30725 17724 30726
rect 17589 30719 17724 30725
rect 17589 30685 17601 30719
rect 17635 30698 17724 30719
rect 17635 30685 17647 30698
rect 17589 30679 17647 30685
rect 14608 30620 15576 30648
rect 14608 30608 14614 30620
rect 16206 30608 16212 30660
rect 16264 30648 16270 30660
rect 16669 30651 16727 30657
rect 16264 30620 16436 30648
rect 16264 30608 16270 30620
rect 14277 30583 14335 30589
rect 14277 30549 14289 30583
rect 14323 30549 14335 30583
rect 14277 30543 14335 30549
rect 14366 30540 14372 30592
rect 14424 30580 14430 30592
rect 16117 30583 16175 30589
rect 16117 30580 16129 30583
rect 14424 30552 16129 30580
rect 14424 30540 14430 30552
rect 16117 30549 16129 30552
rect 16163 30549 16175 30583
rect 16298 30580 16304 30592
rect 16259 30552 16304 30580
rect 16117 30543 16175 30549
rect 16298 30540 16304 30552
rect 16356 30540 16362 30592
rect 16408 30589 16436 30620
rect 16669 30617 16681 30651
rect 16715 30648 16727 30651
rect 16758 30648 16764 30660
rect 16715 30620 16764 30648
rect 16715 30617 16727 30620
rect 16669 30611 16727 30617
rect 16758 30608 16764 30620
rect 16816 30648 16822 30660
rect 17696 30648 17724 30698
rect 19058 30676 19064 30728
rect 19116 30716 19122 30728
rect 19429 30719 19487 30725
rect 19429 30716 19441 30719
rect 19116 30688 19441 30716
rect 19116 30676 19122 30688
rect 19429 30685 19441 30688
rect 19475 30685 19487 30719
rect 19429 30679 19487 30685
rect 19518 30676 19524 30728
rect 19576 30716 19582 30728
rect 20162 30716 20168 30728
rect 19576 30688 19621 30716
rect 20123 30688 20168 30716
rect 19576 30676 19582 30688
rect 20162 30676 20168 30688
rect 20220 30676 20226 30728
rect 20346 30716 20352 30728
rect 20307 30688 20352 30716
rect 20346 30676 20352 30688
rect 20404 30676 20410 30728
rect 16816 30620 17724 30648
rect 18417 30651 18475 30657
rect 16816 30608 16822 30620
rect 18417 30617 18429 30651
rect 18463 30648 18475 30651
rect 19702 30648 19708 30660
rect 18463 30620 19708 30648
rect 18463 30617 18475 30620
rect 18417 30611 18475 30617
rect 19702 30608 19708 30620
rect 19760 30608 19766 30660
rect 20530 30648 20536 30660
rect 19812 30620 20536 30648
rect 16393 30583 16451 30589
rect 16393 30549 16405 30583
rect 16439 30549 16451 30583
rect 16393 30543 16451 30549
rect 16482 30540 16488 30592
rect 16540 30580 16546 30592
rect 16540 30552 16585 30580
rect 16540 30540 16546 30552
rect 17034 30540 17040 30592
rect 17092 30580 17098 30592
rect 18217 30583 18275 30589
rect 18217 30580 18229 30583
rect 17092 30552 18229 30580
rect 17092 30540 17098 30552
rect 18217 30549 18229 30552
rect 18263 30580 18275 30583
rect 19812 30580 19840 30620
rect 20530 30608 20536 30620
rect 20588 30608 20594 30660
rect 20254 30580 20260 30592
rect 18263 30552 19840 30580
rect 20215 30552 20260 30580
rect 18263 30549 18275 30552
rect 18217 30543 18275 30549
rect 20254 30540 20260 30552
rect 20312 30540 20318 30592
rect 1104 30490 29048 30512
rect 1104 30438 7896 30490
rect 7948 30438 7960 30490
rect 8012 30438 8024 30490
rect 8076 30438 8088 30490
rect 8140 30438 8152 30490
rect 8204 30438 14842 30490
rect 14894 30438 14906 30490
rect 14958 30438 14970 30490
rect 15022 30438 15034 30490
rect 15086 30438 15098 30490
rect 15150 30438 21788 30490
rect 21840 30438 21852 30490
rect 21904 30438 21916 30490
rect 21968 30438 21980 30490
rect 22032 30438 22044 30490
rect 22096 30438 28734 30490
rect 28786 30438 28798 30490
rect 28850 30438 28862 30490
rect 28914 30438 28926 30490
rect 28978 30438 28990 30490
rect 29042 30438 29048 30490
rect 1104 30416 29048 30438
rect 5534 30376 5540 30388
rect 2976 30348 3924 30376
rect 2976 30308 3004 30348
rect 3050 30317 3056 30320
rect 2332 30280 3004 30308
rect 2038 30240 2044 30252
rect 1999 30212 2044 30240
rect 2038 30200 2044 30212
rect 2096 30200 2102 30252
rect 2332 30249 2360 30280
rect 3044 30271 3056 30317
rect 3108 30308 3114 30320
rect 3896 30308 3924 30348
rect 4632 30348 5540 30376
rect 4154 30308 4160 30320
rect 3108 30280 3144 30308
rect 3896 30280 4160 30308
rect 3050 30268 3056 30271
rect 3108 30268 3114 30280
rect 4154 30268 4160 30280
rect 4212 30268 4218 30320
rect 2317 30243 2375 30249
rect 2317 30209 2329 30243
rect 2363 30209 2375 30243
rect 3326 30240 3332 30252
rect 2317 30203 2375 30209
rect 2608 30212 3332 30240
rect 2225 30175 2283 30181
rect 2225 30141 2237 30175
rect 2271 30172 2283 30175
rect 2608 30172 2636 30212
rect 3326 30200 3332 30212
rect 3384 30240 3390 30252
rect 4632 30249 4660 30348
rect 5534 30336 5540 30348
rect 5592 30336 5598 30388
rect 8386 30336 8392 30388
rect 8444 30376 8450 30388
rect 10318 30376 10324 30388
rect 8444 30348 10324 30376
rect 8444 30336 8450 30348
rect 10318 30336 10324 30348
rect 10376 30336 10382 30388
rect 10410 30336 10416 30388
rect 10468 30376 10474 30388
rect 10873 30379 10931 30385
rect 10873 30376 10885 30379
rect 10468 30348 10885 30376
rect 10468 30336 10474 30348
rect 10873 30345 10885 30348
rect 10919 30376 10931 30379
rect 11146 30376 11152 30388
rect 10919 30348 11152 30376
rect 10919 30345 10931 30348
rect 10873 30339 10931 30345
rect 11146 30336 11152 30348
rect 11204 30336 11210 30388
rect 12802 30336 12808 30388
rect 12860 30376 12866 30388
rect 14366 30376 14372 30388
rect 12860 30348 14372 30376
rect 12860 30336 12866 30348
rect 14366 30336 14372 30348
rect 14424 30336 14430 30388
rect 15749 30379 15807 30385
rect 14476 30348 15608 30376
rect 6086 30308 6092 30320
rect 4724 30280 6092 30308
rect 4617 30243 4675 30249
rect 3384 30212 4108 30240
rect 3384 30200 3390 30212
rect 2271 30144 2636 30172
rect 2271 30141 2283 30144
rect 2225 30135 2283 30141
rect 2682 30132 2688 30184
rect 2740 30172 2746 30184
rect 2777 30175 2835 30181
rect 2777 30172 2789 30175
rect 2740 30144 2789 30172
rect 2740 30132 2746 30144
rect 2777 30141 2789 30144
rect 2823 30141 2835 30175
rect 2777 30135 2835 30141
rect 1857 30107 1915 30113
rect 1857 30073 1869 30107
rect 1903 30104 1915 30107
rect 1903 30076 2774 30104
rect 1903 30073 1915 30076
rect 1857 30067 1915 30073
rect 2746 30036 2774 30076
rect 3050 30036 3056 30048
rect 2746 30008 3056 30036
rect 3050 29996 3056 30008
rect 3108 29996 3114 30048
rect 4080 30036 4108 30212
rect 4617 30209 4629 30243
rect 4663 30209 4675 30243
rect 4617 30203 4675 30209
rect 4724 30172 4752 30280
rect 6086 30268 6092 30280
rect 6144 30268 6150 30320
rect 6638 30308 6644 30320
rect 6599 30280 6644 30308
rect 6638 30268 6644 30280
rect 6696 30268 6702 30320
rect 7006 30268 7012 30320
rect 7064 30308 7070 30320
rect 12894 30308 12900 30320
rect 7064 30280 12900 30308
rect 7064 30268 7070 30280
rect 12894 30268 12900 30280
rect 12952 30268 12958 30320
rect 14182 30268 14188 30320
rect 14240 30308 14246 30320
rect 14476 30308 14504 30348
rect 14240 30280 14504 30308
rect 14676 30311 14734 30317
rect 14240 30268 14246 30280
rect 14676 30277 14688 30311
rect 14722 30308 14734 30311
rect 14826 30308 14832 30320
rect 14722 30280 14832 30308
rect 14722 30277 14734 30280
rect 14676 30271 14734 30277
rect 14826 30268 14832 30280
rect 14884 30268 14890 30320
rect 15580 30317 15608 30348
rect 15749 30345 15761 30379
rect 15795 30376 15807 30379
rect 15795 30348 16160 30376
rect 15795 30345 15807 30348
rect 15749 30339 15807 30345
rect 15565 30311 15623 30317
rect 15565 30277 15577 30311
rect 15611 30277 15623 30311
rect 15565 30271 15623 30277
rect 4884 30243 4942 30249
rect 4884 30209 4896 30243
rect 4930 30240 4942 30243
rect 5902 30240 5908 30252
rect 4930 30212 5908 30240
rect 4930 30209 4942 30212
rect 4884 30203 4942 30209
rect 5902 30200 5908 30212
rect 5960 30200 5966 30252
rect 6362 30200 6368 30252
rect 6420 30240 6426 30252
rect 6540 30243 6598 30249
rect 6540 30240 6552 30243
rect 6420 30212 6552 30240
rect 6420 30200 6426 30212
rect 6540 30209 6552 30212
rect 6586 30209 6598 30243
rect 6821 30243 6879 30249
rect 6821 30230 6833 30243
rect 6540 30203 6598 30209
rect 6748 30209 6833 30230
rect 6867 30209 6879 30243
rect 6748 30203 6879 30209
rect 6748 30202 6868 30203
rect 4172 30144 4752 30172
rect 4172 30113 4200 30144
rect 6638 30132 6644 30184
rect 6696 30172 6702 30184
rect 6748 30172 6776 30202
rect 7282 30200 7288 30252
rect 7340 30240 7346 30252
rect 7909 30243 7967 30249
rect 7909 30240 7921 30243
rect 7340 30212 7921 30240
rect 7340 30200 7346 30212
rect 7909 30209 7921 30212
rect 7955 30209 7967 30243
rect 7909 30203 7967 30209
rect 9030 30200 9036 30252
rect 9088 30240 9094 30252
rect 9749 30243 9807 30249
rect 9749 30240 9761 30243
rect 9088 30212 9761 30240
rect 9088 30200 9094 30212
rect 9749 30209 9761 30212
rect 9795 30209 9807 30243
rect 9749 30203 9807 30209
rect 10870 30200 10876 30252
rect 10928 30240 10934 30252
rect 11957 30243 12015 30249
rect 11957 30240 11969 30243
rect 10928 30212 11969 30240
rect 10928 30200 10934 30212
rect 11957 30209 11969 30212
rect 12003 30209 12015 30243
rect 11957 30203 12015 30209
rect 12986 30200 12992 30252
rect 13044 30240 13050 30252
rect 14918 30240 14924 30252
rect 13044 30212 14924 30240
rect 13044 30200 13050 30212
rect 14918 30200 14924 30212
rect 14976 30200 14982 30252
rect 15381 30243 15439 30249
rect 15381 30209 15393 30243
rect 15427 30240 15439 30243
rect 15470 30240 15476 30252
rect 15427 30212 15476 30240
rect 15427 30209 15439 30212
rect 15381 30203 15439 30209
rect 15470 30200 15476 30212
rect 15528 30200 15534 30252
rect 15580 30240 15608 30271
rect 15654 30268 15660 30320
rect 15712 30308 15718 30320
rect 16132 30308 16160 30348
rect 16206 30336 16212 30388
rect 16264 30376 16270 30388
rect 16482 30376 16488 30388
rect 16264 30348 16488 30376
rect 16264 30336 16270 30348
rect 16482 30336 16488 30348
rect 16540 30336 16546 30388
rect 17310 30376 17316 30388
rect 16868 30348 17316 30376
rect 16868 30308 16896 30348
rect 17310 30336 17316 30348
rect 17368 30336 17374 30388
rect 17494 30336 17500 30388
rect 17552 30376 17558 30388
rect 17678 30376 17684 30388
rect 17552 30348 17684 30376
rect 17552 30336 17558 30348
rect 17678 30336 17684 30348
rect 17736 30376 17742 30388
rect 19981 30379 20039 30385
rect 19981 30376 19993 30379
rect 17736 30348 19993 30376
rect 17736 30336 17742 30348
rect 19981 30345 19993 30348
rect 20027 30345 20039 30379
rect 19981 30339 20039 30345
rect 19429 30311 19487 30317
rect 19429 30308 19441 30311
rect 15712 30280 15757 30308
rect 16132 30280 16896 30308
rect 17144 30280 19441 30308
rect 15712 30268 15718 30280
rect 17144 30249 17172 30280
rect 19429 30277 19441 30280
rect 19475 30277 19487 30311
rect 19429 30271 19487 30277
rect 19610 30268 19616 30320
rect 19668 30308 19674 30320
rect 20533 30311 20591 30317
rect 20533 30308 20545 30311
rect 19668 30280 20545 30308
rect 19668 30268 19674 30280
rect 20533 30277 20545 30280
rect 20579 30277 20591 30311
rect 20533 30271 20591 30277
rect 17129 30243 17187 30249
rect 15580 30212 17080 30240
rect 7650 30172 7656 30184
rect 6696 30144 6776 30172
rect 7611 30144 7656 30172
rect 6696 30132 6702 30144
rect 7650 30132 7656 30144
rect 7708 30132 7714 30184
rect 9490 30172 9496 30184
rect 9451 30144 9496 30172
rect 9490 30132 9496 30144
rect 9548 30132 9554 30184
rect 11054 30132 11060 30184
rect 11112 30172 11118 30184
rect 11698 30172 11704 30184
rect 11112 30144 11704 30172
rect 11112 30132 11118 30144
rect 11698 30132 11704 30144
rect 11756 30132 11762 30184
rect 16853 30175 16911 30181
rect 16853 30172 16865 30175
rect 15028 30144 16865 30172
rect 4157 30107 4215 30113
rect 4157 30073 4169 30107
rect 4203 30073 4215 30107
rect 4157 30067 4215 30073
rect 5997 30107 6055 30113
rect 5997 30073 6009 30107
rect 6043 30104 6055 30107
rect 6043 30076 7696 30104
rect 6043 30073 6055 30076
rect 5997 30067 6055 30073
rect 6362 30036 6368 30048
rect 4080 30008 6368 30036
rect 6362 29996 6368 30008
rect 6420 29996 6426 30048
rect 6822 30036 6828 30048
rect 6783 30008 6828 30036
rect 6822 29996 6828 30008
rect 6880 29996 6886 30048
rect 7668 30036 7696 30076
rect 13004 30076 13584 30104
rect 8938 30036 8944 30048
rect 7668 30008 8944 30036
rect 8938 29996 8944 30008
rect 8996 29996 9002 30048
rect 9033 30039 9091 30045
rect 9033 30005 9045 30039
rect 9079 30036 9091 30039
rect 10686 30036 10692 30048
rect 9079 30008 10692 30036
rect 9079 30005 9091 30008
rect 9033 29999 9091 30005
rect 10686 29996 10692 30008
rect 10744 29996 10750 30048
rect 10962 29996 10968 30048
rect 11020 30036 11026 30048
rect 13004 30036 13032 30076
rect 11020 30008 13032 30036
rect 11020 29996 11026 30008
rect 13078 29996 13084 30048
rect 13136 30036 13142 30048
rect 13556 30045 13584 30076
rect 13541 30039 13599 30045
rect 13136 30008 13181 30036
rect 13136 29996 13142 30008
rect 13541 30005 13553 30039
rect 13587 30036 13599 30039
rect 15028 30036 15056 30144
rect 16853 30141 16865 30144
rect 16899 30141 16911 30175
rect 17052 30172 17080 30212
rect 17129 30209 17141 30243
rect 17175 30209 17187 30243
rect 17129 30203 17187 30209
rect 17862 30200 17868 30252
rect 17920 30240 17926 30252
rect 17957 30243 18015 30249
rect 17957 30240 17969 30243
rect 17920 30212 17969 30240
rect 17920 30200 17926 30212
rect 17957 30209 17969 30212
rect 18003 30209 18015 30243
rect 17957 30203 18015 30209
rect 18046 30200 18052 30252
rect 18104 30238 18110 30252
rect 18601 30243 18659 30249
rect 18601 30240 18613 30243
rect 18156 30238 18613 30240
rect 18104 30212 18613 30238
rect 18104 30210 18184 30212
rect 18104 30200 18110 30210
rect 18601 30209 18613 30212
rect 18647 30209 18659 30243
rect 18601 30203 18659 30209
rect 19337 30243 19395 30249
rect 19337 30209 19349 30243
rect 19383 30209 19395 30243
rect 19518 30240 19524 30252
rect 19479 30212 19524 30240
rect 19337 30203 19395 30209
rect 17586 30172 17592 30184
rect 17052 30144 17592 30172
rect 16853 30135 16911 30141
rect 17586 30132 17592 30144
rect 17644 30132 17650 30184
rect 18141 30175 18199 30181
rect 18141 30141 18153 30175
rect 18187 30141 18199 30175
rect 18141 30135 18199 30141
rect 15102 30064 15108 30116
rect 15160 30104 15166 30116
rect 15654 30104 15660 30116
rect 15160 30076 15660 30104
rect 15160 30064 15166 30076
rect 15654 30064 15660 30076
rect 15712 30104 15718 30116
rect 17218 30104 17224 30116
rect 15712 30076 17224 30104
rect 15712 30064 15718 30076
rect 17218 30064 17224 30076
rect 17276 30064 17282 30116
rect 13587 30008 15056 30036
rect 13587 30005 13599 30008
rect 13541 29999 13599 30005
rect 15194 29996 15200 30048
rect 15252 30036 15258 30048
rect 15933 30039 15991 30045
rect 15933 30036 15945 30039
rect 15252 30008 15945 30036
rect 15252 29996 15258 30008
rect 15933 30005 15945 30008
rect 15979 30005 15991 30039
rect 16942 30036 16948 30048
rect 16903 30008 16948 30036
rect 15933 29999 15991 30005
rect 16942 29996 16948 30008
rect 17000 29996 17006 30048
rect 17126 29996 17132 30048
rect 17184 30036 17190 30048
rect 17313 30039 17371 30045
rect 17313 30036 17325 30039
rect 17184 30008 17325 30036
rect 17184 29996 17190 30008
rect 17313 30005 17325 30008
rect 17359 30005 17371 30039
rect 17313 29999 17371 30005
rect 17494 29996 17500 30048
rect 17552 30036 17558 30048
rect 17773 30039 17831 30045
rect 17773 30036 17785 30039
rect 17552 30008 17785 30036
rect 17552 29996 17558 30008
rect 17773 30005 17785 30008
rect 17819 30005 17831 30039
rect 17773 29999 17831 30005
rect 18046 29996 18052 30048
rect 18104 30036 18110 30048
rect 18156 30036 18184 30135
rect 18230 30064 18236 30116
rect 18288 30104 18294 30116
rect 18785 30107 18843 30113
rect 18785 30104 18797 30107
rect 18288 30076 18797 30104
rect 18288 30064 18294 30076
rect 18785 30073 18797 30076
rect 18831 30073 18843 30107
rect 18785 30067 18843 30073
rect 18104 30008 18184 30036
rect 18104 29996 18110 30008
rect 18966 29996 18972 30048
rect 19024 30036 19030 30048
rect 19352 30036 19380 30203
rect 19518 30200 19524 30212
rect 19576 30200 19582 30252
rect 28350 30036 28356 30048
rect 19024 30008 19380 30036
rect 28311 30008 28356 30036
rect 19024 29996 19030 30008
rect 28350 29996 28356 30008
rect 28408 29996 28414 30048
rect 1104 29946 28888 29968
rect 1104 29894 4423 29946
rect 4475 29894 4487 29946
rect 4539 29894 4551 29946
rect 4603 29894 4615 29946
rect 4667 29894 4679 29946
rect 4731 29894 11369 29946
rect 11421 29894 11433 29946
rect 11485 29894 11497 29946
rect 11549 29894 11561 29946
rect 11613 29894 11625 29946
rect 11677 29894 18315 29946
rect 18367 29894 18379 29946
rect 18431 29894 18443 29946
rect 18495 29894 18507 29946
rect 18559 29894 18571 29946
rect 18623 29894 25261 29946
rect 25313 29894 25325 29946
rect 25377 29894 25389 29946
rect 25441 29894 25453 29946
rect 25505 29894 25517 29946
rect 25569 29894 28888 29946
rect 1104 29872 28888 29894
rect 6086 29832 6092 29844
rect 4908 29804 6092 29832
rect 3970 29724 3976 29776
rect 4028 29764 4034 29776
rect 4798 29764 4804 29776
rect 4028 29736 4804 29764
rect 4028 29724 4034 29736
rect 4798 29724 4804 29736
rect 4856 29724 4862 29776
rect 4908 29773 4936 29804
rect 6086 29792 6092 29804
rect 6144 29792 6150 29844
rect 6822 29792 6828 29844
rect 6880 29832 6886 29844
rect 9674 29832 9680 29844
rect 6880 29804 9680 29832
rect 6880 29792 6886 29804
rect 9674 29792 9680 29804
rect 9732 29792 9738 29844
rect 13814 29792 13820 29844
rect 13872 29832 13878 29844
rect 13872 29804 14697 29832
rect 13872 29792 13878 29804
rect 4893 29767 4951 29773
rect 4893 29733 4905 29767
rect 4939 29733 4951 29767
rect 4893 29727 4951 29733
rect 6730 29724 6736 29776
rect 6788 29764 6794 29776
rect 7006 29764 7012 29776
rect 6788 29736 7012 29764
rect 6788 29724 6794 29736
rect 7006 29724 7012 29736
rect 7064 29724 7070 29776
rect 7190 29764 7196 29776
rect 7151 29736 7196 29764
rect 7190 29724 7196 29736
rect 7248 29724 7254 29776
rect 10502 29724 10508 29776
rect 10560 29764 10566 29776
rect 11701 29767 11759 29773
rect 10560 29736 11284 29764
rect 10560 29724 10566 29736
rect 5718 29696 5724 29708
rect 4356 29668 5724 29696
rect 2041 29631 2099 29637
rect 2041 29597 2053 29631
rect 2087 29628 2099 29631
rect 2682 29628 2688 29640
rect 2087 29600 2688 29628
rect 2087 29597 2099 29600
rect 2041 29591 2099 29597
rect 2682 29588 2688 29600
rect 2740 29588 2746 29640
rect 2308 29563 2366 29569
rect 2308 29529 2320 29563
rect 2354 29560 2366 29563
rect 2590 29560 2596 29572
rect 2354 29532 2596 29560
rect 2354 29529 2366 29532
rect 2308 29523 2366 29529
rect 2590 29520 2596 29532
rect 2648 29520 2654 29572
rect 4356 29569 4384 29668
rect 5718 29656 5724 29668
rect 5776 29656 5782 29708
rect 6822 29656 6828 29708
rect 6880 29696 6886 29708
rect 7282 29696 7288 29708
rect 6880 29668 7288 29696
rect 6880 29656 6886 29668
rect 7282 29656 7288 29668
rect 7340 29656 7346 29708
rect 10686 29656 10692 29708
rect 10744 29696 10750 29708
rect 10744 29668 11192 29696
rect 10744 29656 10750 29668
rect 4525 29631 4583 29637
rect 4525 29597 4537 29631
rect 4571 29628 4583 29631
rect 5166 29628 5172 29640
rect 4571 29600 5172 29628
rect 4571 29597 4583 29600
rect 4525 29591 4583 29597
rect 5166 29588 5172 29600
rect 5224 29588 5230 29640
rect 6733 29631 6791 29637
rect 6733 29597 6745 29631
rect 6779 29628 6791 29631
rect 8478 29628 8484 29640
rect 6779 29600 8484 29628
rect 6779 29597 6791 29600
rect 6733 29591 6791 29597
rect 8478 29588 8484 29600
rect 8536 29628 8542 29640
rect 8573 29631 8631 29637
rect 8573 29628 8585 29631
rect 8536 29600 8585 29628
rect 8536 29588 8542 29600
rect 8573 29597 8585 29600
rect 8619 29628 8631 29631
rect 9401 29631 9459 29637
rect 9401 29628 9413 29631
rect 8619 29600 9413 29628
rect 8619 29597 8631 29600
rect 8573 29591 8631 29597
rect 9401 29597 9413 29600
rect 9447 29628 9459 29631
rect 9490 29628 9496 29640
rect 9447 29600 9496 29628
rect 9447 29597 9459 29600
rect 9401 29591 9459 29597
rect 9490 29588 9496 29600
rect 9548 29588 9554 29640
rect 10226 29628 10232 29640
rect 9600 29600 10232 29628
rect 4341 29563 4399 29569
rect 4341 29560 4353 29563
rect 2746 29532 4353 29560
rect 1946 29452 1952 29504
rect 2004 29492 2010 29504
rect 2746 29492 2774 29532
rect 4341 29529 4353 29532
rect 4387 29529 4399 29563
rect 4709 29563 4767 29569
rect 4709 29560 4721 29563
rect 4341 29523 4399 29529
rect 4540 29532 4721 29560
rect 2004 29464 2774 29492
rect 3421 29495 3479 29501
rect 2004 29452 2010 29464
rect 3421 29461 3433 29495
rect 3467 29492 3479 29495
rect 3694 29492 3700 29504
rect 3467 29464 3700 29492
rect 3467 29461 3479 29464
rect 3421 29455 3479 29461
rect 3694 29452 3700 29464
rect 3752 29452 3758 29504
rect 4062 29452 4068 29504
rect 4120 29492 4126 29504
rect 4540 29492 4568 29532
rect 4709 29529 4721 29532
rect 4755 29529 4767 29563
rect 6270 29560 6276 29572
rect 4709 29523 4767 29529
rect 5276 29532 6276 29560
rect 4120 29464 4568 29492
rect 4617 29495 4675 29501
rect 4120 29452 4126 29464
rect 4617 29461 4629 29495
rect 4663 29492 4675 29495
rect 5276 29492 5304 29532
rect 6270 29520 6276 29532
rect 6328 29520 6334 29572
rect 6488 29563 6546 29569
rect 6488 29529 6500 29563
rect 6534 29560 6546 29563
rect 7374 29560 7380 29572
rect 6534 29532 7380 29560
rect 6534 29529 6546 29532
rect 6488 29523 6546 29529
rect 7374 29520 7380 29532
rect 7432 29520 7438 29572
rect 8328 29563 8386 29569
rect 8328 29529 8340 29563
rect 8374 29560 8386 29563
rect 9600 29560 9628 29600
rect 10226 29588 10232 29600
rect 10284 29588 10290 29640
rect 10962 29628 10968 29640
rect 10520 29600 10968 29628
rect 8374 29532 9628 29560
rect 9668 29563 9726 29569
rect 8374 29529 8386 29532
rect 8328 29523 8386 29529
rect 9668 29529 9680 29563
rect 9714 29560 9726 29563
rect 9766 29560 9772 29572
rect 9714 29532 9772 29560
rect 9714 29529 9726 29532
rect 9668 29523 9726 29529
rect 9766 29520 9772 29532
rect 9824 29520 9830 29572
rect 4663 29464 5304 29492
rect 5353 29495 5411 29501
rect 4663 29461 4675 29464
rect 4617 29455 4675 29461
rect 5353 29461 5365 29495
rect 5399 29492 5411 29495
rect 7742 29492 7748 29504
rect 5399 29464 7748 29492
rect 5399 29461 5411 29464
rect 5353 29455 5411 29461
rect 7742 29452 7748 29464
rect 7800 29452 7806 29504
rect 8570 29452 8576 29504
rect 8628 29492 8634 29504
rect 10520 29492 10548 29600
rect 10962 29588 10968 29600
rect 11020 29588 11026 29640
rect 10778 29492 10784 29504
rect 8628 29464 10548 29492
rect 10739 29464 10784 29492
rect 8628 29452 8634 29464
rect 10778 29452 10784 29464
rect 10836 29452 10842 29504
rect 11164 29492 11192 29668
rect 11256 29560 11284 29736
rect 11701 29733 11713 29767
rect 11747 29764 11759 29767
rect 11790 29764 11796 29776
rect 11747 29736 11796 29764
rect 11747 29733 11759 29736
rect 11701 29727 11759 29733
rect 11790 29724 11796 29736
rect 11848 29724 11854 29776
rect 13262 29724 13268 29776
rect 13320 29764 13326 29776
rect 13633 29767 13691 29773
rect 13633 29764 13645 29767
rect 13320 29736 13645 29764
rect 13320 29724 13326 29736
rect 13633 29733 13645 29736
rect 13679 29733 13691 29767
rect 14458 29764 14464 29776
rect 13633 29727 13691 29733
rect 14384 29736 14464 29764
rect 13078 29696 13084 29708
rect 13039 29668 13084 29696
rect 13078 29656 13084 29668
rect 13136 29656 13142 29708
rect 11974 29588 11980 29640
rect 12032 29628 12038 29640
rect 14277 29631 14335 29637
rect 14277 29628 14289 29631
rect 12032 29600 14289 29628
rect 12032 29588 12038 29600
rect 14277 29597 14289 29600
rect 14323 29597 14335 29631
rect 14384 29628 14412 29736
rect 14458 29724 14464 29736
rect 14516 29724 14522 29776
rect 14669 29764 14697 29804
rect 14734 29792 14740 29844
rect 14792 29832 14798 29844
rect 15286 29832 15292 29844
rect 14792 29804 15148 29832
rect 15247 29804 15292 29832
rect 14792 29792 14798 29804
rect 15120 29764 15148 29804
rect 15286 29792 15292 29804
rect 15344 29792 15350 29844
rect 15378 29792 15384 29844
rect 15436 29832 15442 29844
rect 15746 29832 15752 29844
rect 15436 29804 15752 29832
rect 15436 29792 15442 29804
rect 15746 29792 15752 29804
rect 15804 29792 15810 29844
rect 17218 29792 17224 29844
rect 17276 29832 17282 29844
rect 17313 29835 17371 29841
rect 17313 29832 17325 29835
rect 17276 29804 17325 29832
rect 17276 29792 17282 29804
rect 17313 29801 17325 29804
rect 17359 29801 17371 29835
rect 20254 29832 20260 29844
rect 17313 29795 17371 29801
rect 17420 29804 18276 29832
rect 15657 29767 15715 29773
rect 14669 29736 14872 29764
rect 15120 29736 15332 29764
rect 14844 29705 14872 29736
rect 15304 29708 15332 29736
rect 15657 29733 15669 29767
rect 15703 29764 15715 29767
rect 15838 29764 15844 29776
rect 15703 29736 15844 29764
rect 15703 29733 15715 29736
rect 15657 29727 15715 29733
rect 15838 29724 15844 29736
rect 15896 29724 15902 29776
rect 15930 29724 15936 29776
rect 15988 29764 15994 29776
rect 17420 29764 17448 29804
rect 15988 29736 17448 29764
rect 15988 29724 15994 29736
rect 17862 29724 17868 29776
rect 17920 29764 17926 29776
rect 18138 29764 18144 29776
rect 17920 29736 18144 29764
rect 17920 29724 17926 29736
rect 18138 29724 18144 29736
rect 18196 29724 18202 29776
rect 18248 29773 18276 29804
rect 19306 29804 20260 29832
rect 18233 29767 18291 29773
rect 18233 29733 18245 29767
rect 18279 29733 18291 29767
rect 18690 29764 18696 29776
rect 18651 29736 18696 29764
rect 18233 29727 18291 29733
rect 18690 29724 18696 29736
rect 18748 29724 18754 29776
rect 14829 29699 14887 29705
rect 14829 29665 14841 29699
rect 14875 29665 14887 29699
rect 14829 29659 14887 29665
rect 14918 29656 14924 29708
rect 14976 29696 14982 29708
rect 15102 29696 15108 29708
rect 14976 29668 15108 29696
rect 14976 29656 14982 29668
rect 15102 29656 15108 29668
rect 15160 29656 15166 29708
rect 15194 29656 15200 29708
rect 15252 29656 15258 29708
rect 15286 29656 15292 29708
rect 15344 29656 15350 29708
rect 15378 29656 15384 29708
rect 15436 29656 15442 29708
rect 19306 29696 19334 29804
rect 20254 29792 20260 29804
rect 20312 29792 20318 29844
rect 16408 29668 19334 29696
rect 14461 29631 14519 29637
rect 14461 29628 14473 29631
rect 14384 29600 14473 29628
rect 14277 29591 14335 29597
rect 14461 29597 14473 29600
rect 14507 29597 14519 29631
rect 14461 29591 14519 29597
rect 14550 29588 14556 29640
rect 14608 29628 14614 29640
rect 14608 29600 14653 29628
rect 14608 29588 14614 29600
rect 14734 29588 14740 29640
rect 14792 29628 14798 29640
rect 15212 29628 15240 29656
rect 14792 29600 15240 29628
rect 15396 29628 15424 29656
rect 15672 29637 15792 29638
rect 15473 29631 15531 29637
rect 15473 29628 15485 29631
rect 15396 29600 15485 29628
rect 14792 29588 14798 29600
rect 15473 29597 15485 29600
rect 15519 29597 15531 29631
rect 15672 29631 15807 29637
rect 15672 29622 15761 29631
rect 15473 29591 15531 29597
rect 15580 29610 15761 29622
rect 15580 29594 15700 29610
rect 15749 29597 15761 29610
rect 15795 29597 15807 29631
rect 16206 29628 16212 29640
rect 16167 29600 16212 29628
rect 12710 29560 12716 29572
rect 11256 29532 12716 29560
rect 12710 29520 12716 29532
rect 12768 29520 12774 29572
rect 12836 29563 12894 29569
rect 12836 29529 12848 29563
rect 12882 29560 12894 29563
rect 13906 29560 13912 29572
rect 12882 29532 13912 29560
rect 12882 29529 12894 29532
rect 12836 29523 12894 29529
rect 13906 29520 13912 29532
rect 13964 29520 13970 29572
rect 15286 29520 15292 29572
rect 15344 29560 15350 29572
rect 15580 29560 15608 29594
rect 15749 29591 15807 29597
rect 16206 29588 16212 29600
rect 16264 29588 16270 29640
rect 16408 29637 16436 29668
rect 16393 29631 16451 29637
rect 16393 29597 16405 29631
rect 16439 29597 16451 29631
rect 16574 29628 16580 29640
rect 16535 29600 16580 29628
rect 16393 29591 16451 29597
rect 16574 29588 16580 29600
rect 16632 29588 16638 29640
rect 16666 29588 16672 29640
rect 16724 29628 16730 29640
rect 16724 29600 16769 29628
rect 16724 29588 16730 29600
rect 17218 29588 17224 29640
rect 17276 29628 17282 29640
rect 17957 29631 18015 29637
rect 17957 29628 17969 29631
rect 17276 29600 17969 29628
rect 17276 29588 17282 29600
rect 17957 29597 17969 29600
rect 18003 29597 18015 29631
rect 18690 29628 18696 29640
rect 18651 29600 18696 29628
rect 17957 29591 18015 29597
rect 18690 29588 18696 29600
rect 18748 29588 18754 29640
rect 18874 29628 18880 29640
rect 18835 29600 18880 29628
rect 18874 29588 18880 29600
rect 18932 29588 18938 29640
rect 28350 29628 28356 29640
rect 28311 29600 28356 29628
rect 28350 29588 28356 29600
rect 28408 29588 28414 29640
rect 15344 29532 15608 29560
rect 15344 29520 15350 29532
rect 16022 29520 16028 29572
rect 16080 29560 16086 29572
rect 17497 29563 17555 29569
rect 16080 29532 17340 29560
rect 16080 29520 16086 29532
rect 17312 29504 17340 29532
rect 17497 29529 17509 29563
rect 17543 29560 17555 29563
rect 17586 29560 17592 29572
rect 17543 29532 17592 29560
rect 17543 29529 17555 29532
rect 17497 29523 17555 29529
rect 17586 29520 17592 29532
rect 17644 29520 17650 29572
rect 17770 29520 17776 29572
rect 17828 29560 17834 29572
rect 18233 29563 18291 29569
rect 18233 29560 18245 29563
rect 17828 29532 18245 29560
rect 17828 29520 17834 29532
rect 18233 29529 18245 29532
rect 18279 29560 18291 29563
rect 19429 29563 19487 29569
rect 19429 29560 19441 29563
rect 18279 29532 19441 29560
rect 18279 29529 18291 29532
rect 18233 29523 18291 29529
rect 19429 29529 19441 29532
rect 19475 29560 19487 29563
rect 19518 29560 19524 29572
rect 19475 29532 19524 29560
rect 19475 29529 19487 29532
rect 19429 29523 19487 29529
rect 19518 29520 19524 29532
rect 19576 29560 19582 29572
rect 19981 29563 20039 29569
rect 19981 29560 19993 29563
rect 19576 29532 19993 29560
rect 19576 29520 19582 29532
rect 19981 29529 19993 29532
rect 20027 29560 20039 29563
rect 20346 29560 20352 29572
rect 20027 29532 20352 29560
rect 20027 29529 20039 29532
rect 19981 29523 20039 29529
rect 20346 29520 20352 29532
rect 20404 29560 20410 29572
rect 20533 29563 20591 29569
rect 20533 29560 20545 29563
rect 20404 29532 20545 29560
rect 20404 29520 20410 29532
rect 20533 29529 20545 29532
rect 20579 29529 20591 29563
rect 20533 29523 20591 29529
rect 13538 29492 13544 29504
rect 11164 29464 13544 29492
rect 13538 29452 13544 29464
rect 13596 29452 13602 29504
rect 14642 29452 14648 29504
rect 14700 29492 14706 29504
rect 17126 29492 17132 29504
rect 14700 29464 14745 29492
rect 17087 29464 17132 29492
rect 14700 29452 14706 29464
rect 17126 29452 17132 29464
rect 17184 29452 17190 29504
rect 17310 29501 17316 29504
rect 17297 29495 17316 29501
rect 17297 29461 17309 29495
rect 17297 29455 17316 29461
rect 17310 29452 17316 29455
rect 17368 29452 17374 29504
rect 18046 29492 18052 29504
rect 18007 29464 18052 29492
rect 18046 29452 18052 29464
rect 18104 29452 18110 29504
rect 1104 29402 29048 29424
rect 1104 29350 7896 29402
rect 7948 29350 7960 29402
rect 8012 29350 8024 29402
rect 8076 29350 8088 29402
rect 8140 29350 8152 29402
rect 8204 29350 14842 29402
rect 14894 29350 14906 29402
rect 14958 29350 14970 29402
rect 15022 29350 15034 29402
rect 15086 29350 15098 29402
rect 15150 29350 21788 29402
rect 21840 29350 21852 29402
rect 21904 29350 21916 29402
rect 21968 29350 21980 29402
rect 22032 29350 22044 29402
rect 22096 29350 28734 29402
rect 28786 29350 28798 29402
rect 28850 29350 28862 29402
rect 28914 29350 28926 29402
rect 28978 29350 28990 29402
rect 29042 29350 29048 29402
rect 1104 29328 29048 29350
rect 2314 29288 2320 29300
rect 2275 29260 2320 29288
rect 2314 29248 2320 29260
rect 2372 29248 2378 29300
rect 3418 29248 3424 29300
rect 3476 29288 3482 29300
rect 5994 29288 6000 29300
rect 3476 29260 5580 29288
rect 5955 29260 6000 29288
rect 3476 29248 3482 29260
rect 2682 29180 2688 29232
rect 2740 29220 2746 29232
rect 5442 29220 5448 29232
rect 2740 29192 5448 29220
rect 2740 29180 2746 29192
rect 1946 29152 1952 29164
rect 1907 29124 1952 29152
rect 1946 29112 1952 29124
rect 2004 29112 2010 29164
rect 2130 29152 2136 29164
rect 2091 29124 2136 29152
rect 2130 29112 2136 29124
rect 2188 29112 2194 29164
rect 2792 29161 2820 29192
rect 3050 29161 3056 29164
rect 2777 29155 2835 29161
rect 2777 29121 2789 29155
rect 2823 29152 2835 29155
rect 2823 29124 2857 29152
rect 2823 29121 2835 29124
rect 2777 29115 2835 29121
rect 3044 29115 3056 29161
rect 3108 29152 3114 29164
rect 4632 29161 4660 29192
rect 5442 29180 5448 29192
rect 5500 29180 5506 29232
rect 5552 29220 5580 29260
rect 5994 29248 6000 29260
rect 6052 29248 6058 29300
rect 6454 29248 6460 29300
rect 6512 29288 6518 29300
rect 7282 29288 7288 29300
rect 6512 29260 7288 29288
rect 6512 29248 6518 29260
rect 7282 29248 7288 29260
rect 7340 29248 7346 29300
rect 7650 29248 7656 29300
rect 7708 29288 7714 29300
rect 8297 29291 8355 29297
rect 8297 29288 8309 29291
rect 7708 29260 8309 29288
rect 7708 29248 7714 29260
rect 8297 29257 8309 29260
rect 8343 29288 8355 29291
rect 11698 29288 11704 29300
rect 8343 29260 11704 29288
rect 8343 29257 8355 29260
rect 8297 29251 8355 29257
rect 11698 29248 11704 29260
rect 11756 29248 11762 29300
rect 11793 29291 11851 29297
rect 11793 29257 11805 29291
rect 11839 29288 11851 29291
rect 12158 29288 12164 29300
rect 11839 29260 12164 29288
rect 11839 29257 11851 29260
rect 11793 29251 11851 29257
rect 12158 29248 12164 29260
rect 12216 29248 12222 29300
rect 12250 29248 12256 29300
rect 12308 29248 12314 29300
rect 12437 29291 12495 29297
rect 12437 29257 12449 29291
rect 12483 29288 12495 29291
rect 12526 29288 12532 29300
rect 12483 29260 12532 29288
rect 12483 29257 12495 29260
rect 12437 29251 12495 29257
rect 12526 29248 12532 29260
rect 12584 29248 12590 29300
rect 12894 29248 12900 29300
rect 12952 29288 12958 29300
rect 14458 29288 14464 29300
rect 12952 29260 14464 29288
rect 12952 29248 12958 29260
rect 14458 29248 14464 29260
rect 14516 29288 14522 29300
rect 14516 29260 14596 29288
rect 14516 29248 14522 29260
rect 9766 29220 9772 29232
rect 5552 29192 9772 29220
rect 9766 29180 9772 29192
rect 9824 29180 9830 29232
rect 11054 29180 11060 29232
rect 11112 29220 11118 29232
rect 12066 29220 12072 29232
rect 11112 29192 12072 29220
rect 11112 29180 11118 29192
rect 12066 29180 12072 29192
rect 12124 29180 12130 29232
rect 12268 29220 12296 29248
rect 12618 29220 12624 29232
rect 12268 29192 12624 29220
rect 12618 29180 12624 29192
rect 12676 29180 12682 29232
rect 14568 29186 14596 29260
rect 14826 29248 14832 29300
rect 14884 29288 14890 29300
rect 15378 29288 15384 29300
rect 14884 29260 15384 29288
rect 14884 29248 14890 29260
rect 15378 29248 15384 29260
rect 15436 29248 15442 29300
rect 16025 29291 16083 29297
rect 16025 29257 16037 29291
rect 16071 29288 16083 29291
rect 16666 29288 16672 29300
rect 16071 29260 16672 29288
rect 16071 29257 16083 29260
rect 16025 29251 16083 29257
rect 16666 29248 16672 29260
rect 16724 29248 16730 29300
rect 17037 29291 17095 29297
rect 17037 29257 17049 29291
rect 17083 29288 17095 29291
rect 18046 29288 18052 29300
rect 17083 29260 18052 29288
rect 17083 29257 17095 29260
rect 17037 29251 17095 29257
rect 14669 29192 15240 29220
rect 14669 29186 14697 29192
rect 4617 29155 4675 29161
rect 3108 29124 3144 29152
rect 3050 29112 3056 29115
rect 3108 29112 3114 29124
rect 4617 29121 4629 29155
rect 4663 29121 4675 29155
rect 4617 29115 4675 29121
rect 4884 29155 4942 29161
rect 4884 29121 4896 29155
rect 4930 29152 4942 29155
rect 5258 29152 5264 29164
rect 4930 29124 5264 29152
rect 4930 29121 4942 29124
rect 4884 29115 4942 29121
rect 5258 29112 5264 29124
rect 5316 29112 5322 29164
rect 5350 29112 5356 29164
rect 5408 29152 5414 29164
rect 5408 29124 6132 29152
rect 5408 29112 5414 29124
rect 1857 29087 1915 29093
rect 1857 29053 1869 29087
rect 1903 29053 1915 29087
rect 1857 29047 1915 29053
rect 1872 29016 1900 29047
rect 4157 29019 4215 29025
rect 1872 28988 2820 29016
rect 4157 28994 4169 29019
rect 2222 28908 2228 28960
rect 2280 28948 2286 28960
rect 2792 28948 2820 28988
rect 4080 28985 4169 28994
rect 4203 28985 4215 29019
rect 6104 29016 6132 29124
rect 6178 29112 6184 29164
rect 6236 29152 6242 29164
rect 6549 29155 6607 29161
rect 6549 29152 6561 29155
rect 6236 29124 6561 29152
rect 6236 29112 6242 29124
rect 6549 29121 6561 29124
rect 6595 29121 6607 29155
rect 6549 29115 6607 29121
rect 7742 29112 7748 29164
rect 7800 29152 7806 29164
rect 8846 29152 8852 29164
rect 7800 29124 8852 29152
rect 7800 29112 7806 29124
rect 8846 29112 8852 29124
rect 8904 29112 8910 29164
rect 9582 29152 9588 29164
rect 9543 29124 9588 29152
rect 9582 29112 9588 29124
rect 9640 29112 9646 29164
rect 9858 29112 9864 29164
rect 9916 29152 9922 29164
rect 10045 29155 10103 29161
rect 10045 29152 10057 29155
rect 9916 29124 10057 29152
rect 9916 29112 9922 29124
rect 10045 29121 10057 29124
rect 10091 29121 10103 29155
rect 10045 29115 10103 29121
rect 11238 29112 11244 29164
rect 11296 29152 11302 29164
rect 12253 29155 12311 29161
rect 12253 29152 12265 29155
rect 11296 29124 12265 29152
rect 11296 29112 11302 29124
rect 12253 29121 12265 29124
rect 12299 29121 12311 29155
rect 12253 29115 12311 29121
rect 12342 29112 12348 29164
rect 12400 29152 12406 29164
rect 12989 29155 13047 29161
rect 14568 29158 14697 29186
rect 12989 29152 13001 29155
rect 12400 29124 13001 29152
rect 12400 29112 12406 29124
rect 12989 29121 13001 29124
rect 13035 29121 13047 29155
rect 12989 29115 13047 29121
rect 14737 29155 14795 29161
rect 14737 29121 14749 29155
rect 14783 29152 14795 29155
rect 15102 29152 15108 29164
rect 14783 29124 15108 29152
rect 14783 29121 14795 29124
rect 14737 29115 14795 29121
rect 15102 29112 15108 29124
rect 15160 29112 15166 29164
rect 15212 29152 15240 29192
rect 15286 29180 15292 29232
rect 15344 29220 15350 29232
rect 17052 29220 17080 29251
rect 18046 29248 18052 29260
rect 18104 29248 18110 29300
rect 15344 29192 17080 29220
rect 15344 29180 15350 29192
rect 15565 29155 15623 29161
rect 15565 29152 15577 29155
rect 15212 29124 15577 29152
rect 15565 29121 15577 29124
rect 15611 29121 15623 29155
rect 15565 29115 15623 29121
rect 15657 29155 15715 29161
rect 15657 29121 15669 29155
rect 15703 29121 15715 29155
rect 15657 29115 15715 29121
rect 15841 29155 15899 29161
rect 15841 29121 15853 29155
rect 15887 29121 15899 29155
rect 16666 29152 16672 29164
rect 15841 29115 15899 29121
rect 16040 29124 16672 29152
rect 6362 29044 6368 29096
rect 6420 29084 6426 29096
rect 6825 29087 6883 29093
rect 6825 29084 6837 29087
rect 6420 29056 6837 29084
rect 6420 29044 6426 29056
rect 6825 29053 6837 29056
rect 6871 29084 6883 29087
rect 7558 29084 7564 29096
rect 6871 29056 7564 29084
rect 6871 29053 6883 29056
rect 6825 29047 6883 29053
rect 7558 29044 7564 29056
rect 7616 29044 7622 29096
rect 11330 29084 11336 29096
rect 7668 29056 11336 29084
rect 7668 29016 7696 29056
rect 11330 29044 11336 29056
rect 11388 29044 11394 29096
rect 11790 29044 11796 29096
rect 11848 29084 11854 29096
rect 14918 29084 14924 29096
rect 11848 29056 14924 29084
rect 11848 29044 11854 29056
rect 14918 29044 14924 29056
rect 14976 29084 14982 29096
rect 15672 29084 15700 29115
rect 14976 29056 15700 29084
rect 14976 29044 14982 29056
rect 6104 28988 7696 29016
rect 4080 28979 4215 28985
rect 4080 28966 4200 28979
rect 7742 28976 7748 29028
rect 7800 29016 7806 29028
rect 8294 29016 8300 29028
rect 7800 28988 8300 29016
rect 7800 28976 7806 28988
rect 8294 28976 8300 28988
rect 8352 28976 8358 29028
rect 8386 28976 8392 29028
rect 8444 29016 8450 29028
rect 10962 29016 10968 29028
rect 8444 28988 10968 29016
rect 8444 28976 8450 28988
rect 10962 28976 10968 28988
rect 11020 28976 11026 29028
rect 11149 29019 11207 29025
rect 11149 28985 11161 29019
rect 11195 29016 11207 29019
rect 12250 29016 12256 29028
rect 11195 28988 12256 29016
rect 11195 28985 11207 28988
rect 11149 28979 11207 28985
rect 12250 28976 12256 28988
rect 12308 28976 12314 29028
rect 15010 29016 15016 29028
rect 12544 28988 15016 29016
rect 2280 28920 2820 28948
rect 2280 28908 2286 28920
rect 3970 28908 3976 28960
rect 4028 28948 4034 28960
rect 4080 28948 4108 28966
rect 4028 28920 4108 28948
rect 4028 28908 4034 28920
rect 10318 28908 10324 28960
rect 10376 28948 10382 28960
rect 11790 28948 11796 28960
rect 10376 28920 11796 28948
rect 10376 28908 10382 28920
rect 11790 28908 11796 28920
rect 11848 28908 11854 28960
rect 11882 28908 11888 28960
rect 11940 28948 11946 28960
rect 12544 28948 12572 28988
rect 15010 28976 15016 28988
rect 15068 28976 15074 29028
rect 15746 29016 15752 29028
rect 15120 28988 15752 29016
rect 11940 28920 12572 28948
rect 11940 28908 11946 28920
rect 12710 28908 12716 28960
rect 12768 28948 12774 28960
rect 15120 28948 15148 28988
rect 15746 28976 15752 28988
rect 15804 28976 15810 29028
rect 15856 29016 15884 29115
rect 16040 29096 16068 29124
rect 16666 29112 16672 29124
rect 16724 29152 16730 29164
rect 16853 29155 16911 29161
rect 16853 29152 16865 29155
rect 16724 29124 16865 29152
rect 16724 29112 16730 29124
rect 16853 29121 16865 29124
rect 16899 29121 16911 29155
rect 16853 29115 16911 29121
rect 17129 29155 17187 29161
rect 17129 29121 17141 29155
rect 17175 29152 17187 29155
rect 17218 29152 17224 29164
rect 17175 29124 17224 29152
rect 17175 29121 17187 29124
rect 17129 29115 17187 29121
rect 16022 29044 16028 29096
rect 16080 29044 16086 29096
rect 16206 29044 16212 29096
rect 16264 29084 16270 29096
rect 17144 29084 17172 29115
rect 17218 29112 17224 29124
rect 17276 29112 17282 29164
rect 17494 29112 17500 29164
rect 17552 29152 17558 29164
rect 17589 29155 17647 29161
rect 17589 29152 17601 29155
rect 17552 29124 17601 29152
rect 17552 29112 17558 29124
rect 17589 29121 17601 29124
rect 17635 29121 17647 29155
rect 17770 29152 17776 29164
rect 17731 29124 17776 29152
rect 17589 29115 17647 29121
rect 17770 29112 17776 29124
rect 17828 29152 17834 29164
rect 18233 29155 18291 29161
rect 18233 29152 18245 29155
rect 17828 29124 18245 29152
rect 17828 29112 17834 29124
rect 18233 29121 18245 29124
rect 18279 29121 18291 29155
rect 18233 29115 18291 29121
rect 16264 29056 17172 29084
rect 16264 29044 16270 29056
rect 16850 29016 16856 29028
rect 15856 28988 16712 29016
rect 16811 28988 16856 29016
rect 12768 28920 15148 28948
rect 12768 28908 12774 28920
rect 15378 28908 15384 28960
rect 15436 28948 15442 28960
rect 16298 28948 16304 28960
rect 15436 28920 16304 28948
rect 15436 28908 15442 28920
rect 16298 28908 16304 28920
rect 16356 28908 16362 28960
rect 16684 28948 16712 28988
rect 16850 28976 16856 28988
rect 16908 28976 16914 29028
rect 17586 29016 17592 29028
rect 17547 28988 17592 29016
rect 17586 28976 17592 28988
rect 17644 28976 17650 29028
rect 18782 29016 18788 29028
rect 17696 28988 18788 29016
rect 17034 28948 17040 28960
rect 16684 28920 17040 28948
rect 17034 28908 17040 28920
rect 17092 28948 17098 28960
rect 17696 28948 17724 28988
rect 18782 28976 18788 28988
rect 18840 28976 18846 29028
rect 17092 28920 17724 28948
rect 17092 28908 17098 28920
rect 1104 28858 28888 28880
rect 1104 28806 4423 28858
rect 4475 28806 4487 28858
rect 4539 28806 4551 28858
rect 4603 28806 4615 28858
rect 4667 28806 4679 28858
rect 4731 28806 11369 28858
rect 11421 28806 11433 28858
rect 11485 28806 11497 28858
rect 11549 28806 11561 28858
rect 11613 28806 11625 28858
rect 11677 28806 18315 28858
rect 18367 28806 18379 28858
rect 18431 28806 18443 28858
rect 18495 28806 18507 28858
rect 18559 28806 18571 28858
rect 18623 28806 25261 28858
rect 25313 28806 25325 28858
rect 25377 28806 25389 28858
rect 25441 28806 25453 28858
rect 25505 28806 25517 28858
rect 25569 28806 28888 28858
rect 1104 28784 28888 28806
rect 5534 28744 5540 28756
rect 5495 28716 5540 28744
rect 5534 28704 5540 28716
rect 5592 28704 5598 28756
rect 6454 28704 6460 28756
rect 6512 28744 6518 28756
rect 8481 28747 8539 28753
rect 8481 28744 8493 28747
rect 6512 28716 8493 28744
rect 6512 28704 6518 28716
rect 8481 28713 8493 28716
rect 8527 28713 8539 28747
rect 8481 28707 8539 28713
rect 9582 28704 9588 28756
rect 9640 28744 9646 28756
rect 11333 28747 11391 28753
rect 11333 28744 11345 28747
rect 9640 28716 11345 28744
rect 9640 28704 9646 28716
rect 11333 28713 11345 28716
rect 11379 28744 11391 28747
rect 12342 28744 12348 28756
rect 11379 28716 12348 28744
rect 11379 28713 11391 28716
rect 11333 28707 11391 28713
rect 12342 28704 12348 28716
rect 12400 28704 12406 28756
rect 13446 28704 13452 28756
rect 13504 28744 13510 28756
rect 13504 28716 14044 28744
rect 13504 28704 13510 28716
rect 3421 28679 3479 28685
rect 3421 28645 3433 28679
rect 3467 28676 3479 28679
rect 6822 28676 6828 28688
rect 3467 28648 6828 28676
rect 3467 28645 3479 28648
rect 3421 28639 3479 28645
rect 6822 28636 6828 28648
rect 6880 28636 6886 28688
rect 8021 28679 8079 28685
rect 8021 28645 8033 28679
rect 8067 28676 8079 28679
rect 8570 28676 8576 28688
rect 8067 28648 8576 28676
rect 8067 28645 8079 28648
rect 8021 28639 8079 28645
rect 8570 28636 8576 28648
rect 8628 28636 8634 28688
rect 9490 28636 9496 28688
rect 9548 28676 9554 28688
rect 9723 28679 9781 28685
rect 9723 28676 9735 28679
rect 9548 28648 9735 28676
rect 9548 28636 9554 28648
rect 9723 28645 9735 28648
rect 9769 28645 9781 28679
rect 12158 28676 12164 28688
rect 9723 28639 9781 28645
rect 9876 28648 12164 28676
rect 9876 28620 9904 28648
rect 12158 28636 12164 28648
rect 12216 28636 12222 28688
rect 12250 28636 12256 28688
rect 12308 28676 12314 28688
rect 14016 28676 14044 28716
rect 14090 28704 14096 28756
rect 14148 28744 14154 28756
rect 14277 28747 14335 28753
rect 14277 28744 14289 28747
rect 14148 28716 14289 28744
rect 14148 28704 14154 28716
rect 14277 28713 14289 28716
rect 14323 28713 14335 28747
rect 14277 28707 14335 28713
rect 15381 28747 15439 28753
rect 15381 28713 15393 28747
rect 15427 28744 15439 28747
rect 15470 28744 15476 28756
rect 15427 28716 15476 28744
rect 15427 28713 15439 28716
rect 15381 28707 15439 28713
rect 15470 28704 15476 28716
rect 15528 28704 15534 28756
rect 15749 28747 15807 28753
rect 15749 28713 15761 28747
rect 15795 28744 15807 28747
rect 16114 28744 16120 28756
rect 15795 28716 16120 28744
rect 15795 28713 15807 28716
rect 15749 28707 15807 28713
rect 16114 28704 16120 28716
rect 16172 28704 16178 28756
rect 16485 28747 16543 28753
rect 16485 28713 16497 28747
rect 16531 28744 16543 28747
rect 18690 28744 18696 28756
rect 16531 28716 18696 28744
rect 16531 28713 16543 28716
rect 16485 28707 16543 28713
rect 18690 28704 18696 28716
rect 18748 28704 18754 28756
rect 12308 28648 13584 28676
rect 14016 28648 15884 28676
rect 12308 28636 12314 28648
rect 7469 28611 7527 28617
rect 7469 28577 7481 28611
rect 7515 28608 7527 28611
rect 9858 28608 9864 28620
rect 7515 28580 9864 28608
rect 7515 28577 7527 28580
rect 7469 28571 7527 28577
rect 9858 28568 9864 28580
rect 9916 28568 9922 28620
rect 9953 28611 10011 28617
rect 9953 28577 9965 28611
rect 9999 28608 10011 28611
rect 13170 28608 13176 28620
rect 9999 28580 13176 28608
rect 9999 28577 10011 28580
rect 9953 28571 10011 28577
rect 13170 28568 13176 28580
rect 13228 28568 13234 28620
rect 2041 28543 2099 28549
rect 2041 28509 2053 28543
rect 2087 28540 2099 28543
rect 2682 28540 2688 28552
rect 2087 28512 2688 28540
rect 2087 28509 2099 28512
rect 2041 28503 2099 28509
rect 2682 28500 2688 28512
rect 2740 28500 2746 28552
rect 4801 28543 4859 28549
rect 4801 28509 4813 28543
rect 4847 28540 4859 28543
rect 5810 28540 5816 28552
rect 4847 28512 5816 28540
rect 4847 28509 4859 28512
rect 4801 28503 4859 28509
rect 5810 28500 5816 28512
rect 5868 28500 5874 28552
rect 7009 28543 7067 28549
rect 7009 28509 7021 28543
rect 7055 28540 7067 28543
rect 9582 28540 9588 28552
rect 7055 28512 9588 28540
rect 7055 28509 7067 28512
rect 7009 28503 7067 28509
rect 9582 28500 9588 28512
rect 9640 28500 9646 28552
rect 9766 28500 9772 28552
rect 9824 28540 9830 28552
rect 13265 28543 13323 28549
rect 13265 28540 13277 28543
rect 9824 28512 13277 28540
rect 9824 28500 9830 28512
rect 13265 28509 13277 28512
rect 13311 28509 13323 28543
rect 13265 28503 13323 28509
rect 13449 28543 13507 28549
rect 13449 28509 13461 28543
rect 13495 28540 13507 28543
rect 13556 28540 13584 28648
rect 13630 28568 13636 28620
rect 13688 28608 13694 28620
rect 13688 28580 13733 28608
rect 13688 28568 13694 28580
rect 14274 28568 14280 28620
rect 14332 28608 14338 28620
rect 14568 28617 14596 28648
rect 14436 28611 14494 28617
rect 14436 28608 14448 28611
rect 14332 28580 14448 28608
rect 14332 28568 14338 28580
rect 14436 28577 14448 28580
rect 14482 28577 14494 28611
rect 14436 28571 14494 28577
rect 14553 28611 14611 28617
rect 14553 28577 14565 28611
rect 14599 28577 14611 28611
rect 14553 28571 14611 28577
rect 14645 28611 14703 28617
rect 14645 28577 14657 28611
rect 14691 28608 14703 28611
rect 14734 28608 14740 28620
rect 14691 28580 14740 28608
rect 14691 28577 14703 28580
rect 14645 28571 14703 28577
rect 14734 28568 14740 28580
rect 14792 28568 14798 28620
rect 14918 28608 14924 28620
rect 14879 28580 14924 28608
rect 14918 28568 14924 28580
rect 14976 28568 14982 28620
rect 15856 28617 15884 28648
rect 16298 28636 16304 28688
rect 16356 28676 16362 28688
rect 17037 28679 17095 28685
rect 17037 28676 17049 28679
rect 16356 28648 17049 28676
rect 16356 28636 16362 28648
rect 17037 28645 17049 28648
rect 17083 28645 17095 28679
rect 17037 28639 17095 28645
rect 18138 28636 18144 28688
rect 18196 28676 18202 28688
rect 18233 28679 18291 28685
rect 18233 28676 18245 28679
rect 18196 28648 18245 28676
rect 18196 28636 18202 28648
rect 18233 28645 18245 28648
rect 18279 28645 18291 28679
rect 18233 28639 18291 28645
rect 15841 28611 15899 28617
rect 15841 28577 15853 28611
rect 15887 28577 15899 28611
rect 15841 28571 15899 28577
rect 15930 28568 15936 28620
rect 15988 28608 15994 28620
rect 16393 28611 16451 28617
rect 16393 28608 16405 28611
rect 15988 28580 16405 28608
rect 15988 28568 15994 28580
rect 16393 28577 16405 28580
rect 16439 28577 16451 28611
rect 16574 28608 16580 28620
rect 16535 28580 16580 28608
rect 16393 28571 16451 28577
rect 16574 28568 16580 28580
rect 16632 28568 16638 28620
rect 13495 28512 13952 28540
rect 13495 28509 13507 28512
rect 13449 28503 13507 28509
rect 2308 28475 2366 28481
rect 2308 28441 2320 28475
rect 2354 28472 2366 28475
rect 4157 28475 4215 28481
rect 4157 28472 4169 28475
rect 2354 28444 4169 28472
rect 2354 28441 2366 28444
rect 2308 28435 2366 28441
rect 4157 28441 4169 28444
rect 4203 28441 4215 28475
rect 4157 28435 4215 28441
rect 4430 28432 4436 28484
rect 4488 28472 4494 28484
rect 5442 28472 5448 28484
rect 4488 28444 5448 28472
rect 4488 28432 4494 28444
rect 5442 28432 5448 28444
rect 5500 28472 5506 28484
rect 7098 28472 7104 28484
rect 5500 28444 7104 28472
rect 5500 28432 5506 28444
rect 7098 28432 7104 28444
rect 7156 28432 7162 28484
rect 7653 28475 7711 28481
rect 7653 28472 7665 28475
rect 7484 28444 7665 28472
rect 4062 28364 4068 28416
rect 4120 28404 4126 28416
rect 7484 28404 7512 28444
rect 7653 28441 7665 28444
rect 7699 28472 7711 28475
rect 8570 28472 8576 28484
rect 7699 28444 8576 28472
rect 7699 28441 7711 28444
rect 7653 28435 7711 28441
rect 8570 28432 8576 28444
rect 8628 28432 8634 28484
rect 8662 28432 8668 28484
rect 8720 28472 8726 28484
rect 12250 28472 12256 28484
rect 8720 28444 12256 28472
rect 8720 28432 8726 28444
rect 12250 28432 12256 28444
rect 12308 28432 12314 28484
rect 12618 28472 12624 28484
rect 12579 28444 12624 28472
rect 12618 28432 12624 28444
rect 12676 28432 12682 28484
rect 13814 28472 13820 28484
rect 13004 28444 13308 28472
rect 4120 28376 7512 28404
rect 4120 28364 4126 28376
rect 7558 28364 7564 28416
rect 7616 28404 7622 28416
rect 7745 28407 7803 28413
rect 7745 28404 7757 28407
rect 7616 28376 7757 28404
rect 7616 28364 7622 28376
rect 7745 28373 7757 28376
rect 7791 28373 7803 28407
rect 7745 28367 7803 28373
rect 7837 28407 7895 28413
rect 7837 28373 7849 28407
rect 7883 28404 7895 28407
rect 10686 28404 10692 28416
rect 7883 28376 10692 28404
rect 7883 28373 7895 28376
rect 7837 28367 7895 28373
rect 10686 28364 10692 28376
rect 10744 28364 10750 28416
rect 10962 28364 10968 28416
rect 11020 28404 11026 28416
rect 12066 28404 12072 28416
rect 11020 28376 12072 28404
rect 11020 28364 11026 28376
rect 12066 28364 12072 28376
rect 12124 28404 12130 28416
rect 13004 28404 13032 28444
rect 12124 28376 13032 28404
rect 13081 28407 13139 28413
rect 12124 28364 12130 28376
rect 13081 28373 13093 28407
rect 13127 28404 13139 28407
rect 13170 28404 13176 28416
rect 13127 28376 13176 28404
rect 13127 28373 13139 28376
rect 13081 28367 13139 28373
rect 13170 28364 13176 28376
rect 13228 28364 13234 28416
rect 13280 28404 13308 28444
rect 13648 28444 13820 28472
rect 13357 28407 13415 28413
rect 13357 28404 13369 28407
rect 13280 28376 13369 28404
rect 13357 28373 13369 28376
rect 13403 28404 13415 28407
rect 13648 28404 13676 28444
rect 13814 28432 13820 28444
rect 13872 28432 13878 28484
rect 13924 28472 13952 28512
rect 13998 28500 14004 28552
rect 14056 28540 14062 28552
rect 15565 28543 15623 28549
rect 15565 28540 15577 28543
rect 14056 28512 15577 28540
rect 14056 28500 14062 28512
rect 15565 28509 15577 28512
rect 15611 28509 15623 28543
rect 15565 28503 15623 28509
rect 16301 28543 16359 28549
rect 16301 28509 16313 28543
rect 16347 28509 16359 28543
rect 16301 28503 16359 28509
rect 14090 28472 14096 28484
rect 13924 28444 14096 28472
rect 14090 28432 14096 28444
rect 14148 28432 14154 28484
rect 14200 28444 14412 28472
rect 13403 28376 13676 28404
rect 13403 28373 13415 28376
rect 13357 28367 13415 28373
rect 13722 28364 13728 28416
rect 13780 28404 13786 28416
rect 14200 28404 14228 28444
rect 13780 28376 14228 28404
rect 14384 28404 14412 28444
rect 14568 28444 15792 28472
rect 14568 28404 14596 28444
rect 14384 28376 14596 28404
rect 15764 28404 15792 28444
rect 15838 28432 15844 28484
rect 15896 28472 15902 28484
rect 16316 28472 16344 28503
rect 16942 28500 16948 28552
rect 17000 28540 17006 28552
rect 17037 28543 17095 28549
rect 17037 28540 17049 28543
rect 17000 28512 17049 28540
rect 17000 28500 17006 28512
rect 17037 28509 17049 28512
rect 17083 28509 17095 28543
rect 17037 28503 17095 28509
rect 17221 28543 17279 28549
rect 17221 28509 17233 28543
rect 17267 28540 17279 28543
rect 17310 28540 17316 28552
rect 17267 28512 17316 28540
rect 17267 28509 17279 28512
rect 17221 28503 17279 28509
rect 15896 28444 16344 28472
rect 15896 28432 15902 28444
rect 17052 28404 17080 28503
rect 17310 28500 17316 28512
rect 17368 28540 17374 28552
rect 17681 28543 17739 28549
rect 17681 28540 17693 28543
rect 17368 28512 17693 28540
rect 17368 28500 17374 28512
rect 17681 28509 17693 28512
rect 17727 28540 17739 28543
rect 17770 28540 17776 28552
rect 17727 28512 17776 28540
rect 17727 28509 17739 28512
rect 17681 28503 17739 28509
rect 17770 28500 17776 28512
rect 17828 28500 17834 28552
rect 15764 28376 17080 28404
rect 13780 28364 13786 28376
rect 1104 28314 29048 28336
rect 1104 28262 7896 28314
rect 7948 28262 7960 28314
rect 8012 28262 8024 28314
rect 8076 28262 8088 28314
rect 8140 28262 8152 28314
rect 8204 28262 14842 28314
rect 14894 28262 14906 28314
rect 14958 28262 14970 28314
rect 15022 28262 15034 28314
rect 15086 28262 15098 28314
rect 15150 28262 21788 28314
rect 21840 28262 21852 28314
rect 21904 28262 21916 28314
rect 21968 28262 21980 28314
rect 22032 28262 22044 28314
rect 22096 28262 28734 28314
rect 28786 28262 28798 28314
rect 28850 28262 28862 28314
rect 28914 28262 28926 28314
rect 28978 28262 28990 28314
rect 29042 28262 29048 28314
rect 1104 28240 29048 28262
rect 5626 28200 5632 28212
rect 3344 28172 5632 28200
rect 3176 28135 3234 28141
rect 3176 28101 3188 28135
rect 3222 28132 3234 28135
rect 3344 28132 3372 28172
rect 5626 28160 5632 28172
rect 5684 28160 5690 28212
rect 5810 28160 5816 28212
rect 5868 28200 5874 28212
rect 8294 28200 8300 28212
rect 5868 28172 8300 28200
rect 5868 28160 5874 28172
rect 8294 28160 8300 28172
rect 8352 28200 8358 28212
rect 8941 28203 8999 28209
rect 8941 28200 8953 28203
rect 8352 28172 8953 28200
rect 8352 28160 8358 28172
rect 8941 28169 8953 28172
rect 8987 28169 8999 28203
rect 8941 28163 8999 28169
rect 10781 28203 10839 28209
rect 10781 28169 10793 28203
rect 10827 28200 10839 28203
rect 12894 28200 12900 28212
rect 10827 28172 12900 28200
rect 10827 28169 10839 28172
rect 10781 28163 10839 28169
rect 12894 28160 12900 28172
rect 12952 28160 12958 28212
rect 12986 28160 12992 28212
rect 13044 28200 13050 28212
rect 13170 28200 13176 28212
rect 13044 28172 13176 28200
rect 13044 28160 13050 28172
rect 13170 28160 13176 28172
rect 13228 28200 13234 28212
rect 15930 28200 15936 28212
rect 13228 28172 15936 28200
rect 13228 28160 13234 28172
rect 15930 28160 15936 28172
rect 15988 28160 15994 28212
rect 5534 28132 5540 28144
rect 3222 28104 3372 28132
rect 3436 28104 5540 28132
rect 3222 28101 3234 28104
rect 3176 28095 3234 28101
rect 3436 28073 3464 28104
rect 3421 28067 3479 28073
rect 3421 28033 3433 28067
rect 3467 28033 3479 28067
rect 3421 28027 3479 28033
rect 4065 28067 4123 28073
rect 4065 28033 4077 28067
rect 4111 28064 4123 28067
rect 4430 28064 4436 28076
rect 4111 28036 4436 28064
rect 4111 28033 4123 28036
rect 4065 28027 4123 28033
rect 4430 28024 4436 28036
rect 4488 28024 4494 28076
rect 4632 28073 4660 28104
rect 5534 28092 5540 28104
rect 5592 28092 5598 28144
rect 8478 28132 8484 28144
rect 7576 28104 8484 28132
rect 4890 28073 4896 28076
rect 4617 28067 4675 28073
rect 4617 28033 4629 28067
rect 4663 28033 4675 28067
rect 4617 28027 4675 28033
rect 4884 28027 4896 28073
rect 4948 28064 4954 28076
rect 4948 28036 4984 28064
rect 4890 28024 4896 28027
rect 4948 28024 4954 28036
rect 5718 28024 5724 28076
rect 5776 28064 5782 28076
rect 6733 28067 6791 28073
rect 6733 28064 6745 28067
rect 5776 28036 6745 28064
rect 5776 28024 5782 28036
rect 6733 28033 6745 28036
rect 6779 28064 6791 28067
rect 7098 28064 7104 28076
rect 6779 28036 7104 28064
rect 6779 28033 6791 28036
rect 6733 28027 6791 28033
rect 7098 28024 7104 28036
rect 7156 28024 7162 28076
rect 7576 28073 7604 28104
rect 8478 28092 8484 28104
rect 8536 28092 8542 28144
rect 9668 28135 9726 28141
rect 9668 28101 9680 28135
rect 9714 28132 9726 28135
rect 9950 28132 9956 28144
rect 9714 28104 9956 28132
rect 9714 28101 9726 28104
rect 9668 28095 9726 28101
rect 9950 28092 9956 28104
rect 10008 28092 10014 28144
rect 14829 28135 14887 28141
rect 14829 28132 14841 28135
rect 12084 28104 14841 28132
rect 7561 28067 7619 28073
rect 7561 28033 7573 28067
rect 7607 28033 7619 28067
rect 7561 28027 7619 28033
rect 7650 28024 7656 28076
rect 7708 28064 7714 28076
rect 7817 28067 7875 28073
rect 7817 28064 7829 28067
rect 7708 28036 7829 28064
rect 7708 28024 7714 28036
rect 7817 28033 7829 28036
rect 7863 28033 7875 28067
rect 8496 28064 8524 28092
rect 9401 28067 9459 28073
rect 9401 28064 9413 28067
rect 8496 28036 9413 28064
rect 7817 28027 7875 28033
rect 9401 28033 9413 28036
rect 9447 28033 9459 28067
rect 9401 28027 9459 28033
rect 11968 28067 12026 28073
rect 11968 28033 11980 28067
rect 12014 28064 12026 28067
rect 12084 28064 12112 28104
rect 14829 28101 14841 28104
rect 14875 28101 14887 28135
rect 14829 28095 14887 28101
rect 12014 28036 12112 28064
rect 14093 28067 14151 28073
rect 12014 28033 12026 28036
rect 11968 28027 12026 28033
rect 14093 28033 14105 28067
rect 14139 28064 14151 28067
rect 14734 28064 14740 28076
rect 14139 28036 14740 28064
rect 14139 28033 14151 28036
rect 14093 28027 14151 28033
rect 14734 28024 14740 28036
rect 14792 28024 14798 28076
rect 15010 28064 15016 28076
rect 14971 28036 15016 28064
rect 15010 28024 15016 28036
rect 15068 28024 15074 28076
rect 15838 28064 15844 28076
rect 15120 28036 15844 28064
rect 6454 27956 6460 28008
rect 6512 27996 6518 28008
rect 6825 27999 6883 28005
rect 6825 27996 6837 27999
rect 6512 27968 6837 27996
rect 6512 27956 6518 27968
rect 6825 27965 6837 27968
rect 6871 27965 6883 27999
rect 6825 27959 6883 27965
rect 6917 27999 6975 28005
rect 6917 27965 6929 27999
rect 6963 27965 6975 27999
rect 6917 27959 6975 27965
rect 7009 27999 7067 28005
rect 7009 27965 7021 27999
rect 7055 27996 7067 27999
rect 7190 27996 7196 28008
rect 7055 27968 7196 27996
rect 7055 27965 7067 27968
rect 7009 27959 7067 27965
rect 3602 27888 3608 27940
rect 3660 27928 3666 27940
rect 3881 27931 3939 27937
rect 3881 27928 3893 27931
rect 3660 27900 3893 27928
rect 3660 27888 3666 27900
rect 3881 27897 3893 27900
rect 3927 27897 3939 27931
rect 6549 27931 6607 27937
rect 6549 27928 6561 27931
rect 3881 27891 3939 27897
rect 5552 27900 6561 27928
rect 2041 27863 2099 27869
rect 2041 27829 2053 27863
rect 2087 27860 2099 27863
rect 2314 27860 2320 27872
rect 2087 27832 2320 27860
rect 2087 27829 2099 27832
rect 2041 27823 2099 27829
rect 2314 27820 2320 27832
rect 2372 27820 2378 27872
rect 4154 27820 4160 27872
rect 4212 27860 4218 27872
rect 5552 27860 5580 27900
rect 6549 27897 6561 27900
rect 6595 27897 6607 27931
rect 6932 27928 6960 27959
rect 7190 27956 7196 27968
rect 7248 27956 7254 28008
rect 11698 27996 11704 28008
rect 11659 27968 11704 27996
rect 11698 27956 11704 27968
rect 11756 27956 11762 28008
rect 14366 27996 14372 28008
rect 14327 27968 14372 27996
rect 14366 27956 14372 27968
rect 14424 27956 14430 28008
rect 15120 27996 15148 28036
rect 15838 28024 15844 28036
rect 15896 28024 15902 28076
rect 15930 28024 15936 28076
rect 15988 28064 15994 28076
rect 15988 28036 16033 28064
rect 15988 28024 15994 28036
rect 14476 27968 15148 27996
rect 15289 27999 15347 28005
rect 7558 27928 7564 27940
rect 6932 27900 7564 27928
rect 6549 27891 6607 27897
rect 7558 27888 7564 27900
rect 7616 27888 7622 27940
rect 12710 27888 12716 27940
rect 12768 27928 12774 27940
rect 14476 27928 14504 27968
rect 15289 27965 15301 27999
rect 15335 27996 15347 27999
rect 15470 27996 15476 28008
rect 15335 27968 15476 27996
rect 15335 27965 15347 27968
rect 15289 27959 15347 27965
rect 15470 27956 15476 27968
rect 15528 27996 15534 28008
rect 16482 27996 16488 28008
rect 15528 27968 16488 27996
rect 15528 27956 15534 27968
rect 16482 27956 16488 27968
rect 16540 27956 16546 28008
rect 12768 27900 14504 27928
rect 12768 27888 12774 27900
rect 15102 27888 15108 27940
rect 15160 27928 15166 27940
rect 16574 27928 16580 27940
rect 15160 27900 16580 27928
rect 15160 27888 15166 27900
rect 16574 27888 16580 27900
rect 16632 27928 16638 27940
rect 16853 27931 16911 27937
rect 16853 27928 16865 27931
rect 16632 27900 16865 27928
rect 16632 27888 16638 27900
rect 16853 27897 16865 27900
rect 16899 27897 16911 27931
rect 16853 27891 16911 27897
rect 4212 27832 5580 27860
rect 5997 27863 6055 27869
rect 4212 27820 4218 27832
rect 5997 27829 6009 27863
rect 6043 27860 6055 27863
rect 6086 27860 6092 27872
rect 6043 27832 6092 27860
rect 6043 27829 6055 27832
rect 5997 27823 6055 27829
rect 6086 27820 6092 27832
rect 6144 27860 6150 27872
rect 6362 27860 6368 27872
rect 6144 27832 6368 27860
rect 6144 27820 6150 27832
rect 6362 27820 6368 27832
rect 6420 27820 6426 27872
rect 8570 27820 8576 27872
rect 8628 27860 8634 27872
rect 12986 27860 12992 27872
rect 8628 27832 12992 27860
rect 8628 27820 8634 27832
rect 12986 27820 12992 27832
rect 13044 27820 13050 27872
rect 13081 27863 13139 27869
rect 13081 27829 13093 27863
rect 13127 27860 13139 27863
rect 13262 27860 13268 27872
rect 13127 27832 13268 27860
rect 13127 27829 13139 27832
rect 13081 27823 13139 27829
rect 13262 27820 13268 27832
rect 13320 27860 13326 27872
rect 13446 27860 13452 27872
rect 13320 27832 13452 27860
rect 13320 27820 13326 27832
rect 13446 27820 13452 27832
rect 13504 27820 13510 27872
rect 13906 27860 13912 27872
rect 13867 27832 13912 27860
rect 13906 27820 13912 27832
rect 13964 27820 13970 27872
rect 14274 27860 14280 27872
rect 14235 27832 14280 27860
rect 14274 27820 14280 27832
rect 14332 27820 14338 27872
rect 15197 27863 15255 27869
rect 15197 27829 15209 27863
rect 15243 27860 15255 27863
rect 15378 27860 15384 27872
rect 15243 27832 15384 27860
rect 15243 27829 15255 27832
rect 15197 27823 15255 27829
rect 15378 27820 15384 27832
rect 15436 27820 15442 27872
rect 16022 27820 16028 27872
rect 16080 27860 16086 27872
rect 16117 27863 16175 27869
rect 16117 27860 16129 27863
rect 16080 27832 16129 27860
rect 16080 27820 16086 27832
rect 16117 27829 16129 27832
rect 16163 27860 16175 27863
rect 18874 27860 18880 27872
rect 16163 27832 18880 27860
rect 16163 27829 16175 27832
rect 16117 27823 16175 27829
rect 18874 27820 18880 27832
rect 18932 27820 18938 27872
rect 28350 27860 28356 27872
rect 28311 27832 28356 27860
rect 28350 27820 28356 27832
rect 28408 27820 28414 27872
rect 1104 27770 28888 27792
rect 1104 27718 4423 27770
rect 4475 27718 4487 27770
rect 4539 27718 4551 27770
rect 4603 27718 4615 27770
rect 4667 27718 4679 27770
rect 4731 27718 11369 27770
rect 11421 27718 11433 27770
rect 11485 27718 11497 27770
rect 11549 27718 11561 27770
rect 11613 27718 11625 27770
rect 11677 27718 18315 27770
rect 18367 27718 18379 27770
rect 18431 27718 18443 27770
rect 18495 27718 18507 27770
rect 18559 27718 18571 27770
rect 18623 27718 25261 27770
rect 25313 27718 25325 27770
rect 25377 27718 25389 27770
rect 25441 27718 25453 27770
rect 25505 27718 25517 27770
rect 25569 27718 28888 27770
rect 1104 27696 28888 27718
rect 4341 27659 4399 27665
rect 4341 27625 4353 27659
rect 4387 27656 4399 27659
rect 4890 27656 4896 27668
rect 4387 27628 4896 27656
rect 4387 27625 4399 27628
rect 4341 27619 4399 27625
rect 4890 27616 4896 27628
rect 4948 27616 4954 27668
rect 6086 27656 6092 27668
rect 5276 27628 6092 27656
rect 3418 27588 3424 27600
rect 3379 27560 3424 27588
rect 3418 27548 3424 27560
rect 3476 27548 3482 27600
rect 5166 27588 5172 27600
rect 4724 27560 5172 27588
rect 1949 27523 2007 27529
rect 1949 27489 1961 27523
rect 1995 27520 2007 27523
rect 2590 27520 2596 27532
rect 1995 27492 2596 27520
rect 1995 27489 2007 27492
rect 1949 27483 2007 27489
rect 2590 27480 2596 27492
rect 2648 27480 2654 27532
rect 4724 27520 4752 27560
rect 5166 27548 5172 27560
rect 5224 27548 5230 27600
rect 2792 27492 4752 27520
rect 4813 27523 4871 27529
rect 2133 27455 2191 27461
rect 2133 27421 2145 27455
rect 2179 27452 2191 27455
rect 2792 27452 2820 27492
rect 4813 27489 4825 27523
rect 4859 27520 4871 27523
rect 5276 27520 5304 27628
rect 6086 27616 6092 27628
rect 6144 27616 6150 27668
rect 7466 27616 7472 27668
rect 7524 27656 7530 27668
rect 12250 27656 12256 27668
rect 7524 27628 12256 27656
rect 7524 27616 7530 27628
rect 12250 27616 12256 27628
rect 12308 27616 12314 27668
rect 12342 27616 12348 27668
rect 12400 27656 12406 27668
rect 15102 27656 15108 27668
rect 12400 27628 15108 27656
rect 12400 27616 12406 27628
rect 15102 27616 15108 27628
rect 15160 27616 15166 27668
rect 15286 27656 15292 27668
rect 15247 27628 15292 27656
rect 15286 27616 15292 27628
rect 15344 27616 15350 27668
rect 5350 27548 5356 27600
rect 5408 27588 5414 27600
rect 11241 27591 11299 27597
rect 5408 27560 5453 27588
rect 5408 27548 5414 27560
rect 11241 27557 11253 27591
rect 11287 27588 11299 27591
rect 11606 27588 11612 27600
rect 11287 27560 11612 27588
rect 11287 27557 11299 27560
rect 11241 27551 11299 27557
rect 11606 27548 11612 27560
rect 11664 27588 11670 27600
rect 11664 27560 11836 27588
rect 11664 27548 11670 27560
rect 5718 27520 5724 27532
rect 4859 27492 5304 27520
rect 5460 27492 5724 27520
rect 4859 27489 4871 27492
rect 4813 27483 4871 27489
rect 3326 27452 3332 27464
rect 2179 27424 2820 27452
rect 3287 27424 3332 27452
rect 2179 27421 2191 27424
rect 2133 27415 2191 27421
rect 3326 27412 3332 27424
rect 3384 27412 3390 27464
rect 3421 27455 3479 27461
rect 3421 27421 3433 27455
rect 3467 27452 3479 27455
rect 4062 27452 4068 27464
rect 3467 27424 4068 27452
rect 3467 27421 3479 27424
rect 3421 27415 3479 27421
rect 4062 27412 4068 27424
rect 4120 27412 4126 27464
rect 4525 27455 4583 27461
rect 4525 27421 4537 27455
rect 4571 27452 4583 27455
rect 4614 27452 4620 27464
rect 4571 27424 4620 27452
rect 4571 27421 4583 27424
rect 4525 27415 4583 27421
rect 4614 27412 4620 27424
rect 4672 27412 4678 27464
rect 4709 27455 4767 27461
rect 4709 27421 4721 27455
rect 4755 27452 4767 27455
rect 5460 27452 5488 27492
rect 5718 27480 5724 27492
rect 5776 27480 5782 27532
rect 10689 27523 10747 27529
rect 10689 27489 10701 27523
rect 10735 27520 10747 27523
rect 11698 27520 11704 27532
rect 10735 27492 11704 27520
rect 10735 27489 10747 27492
rect 10689 27483 10747 27489
rect 11698 27480 11704 27492
rect 11756 27480 11762 27532
rect 11808 27520 11836 27560
rect 11882 27548 11888 27600
rect 11940 27588 11946 27600
rect 14366 27588 14372 27600
rect 11940 27560 14372 27588
rect 11940 27548 11946 27560
rect 14366 27548 14372 27560
rect 14424 27548 14430 27600
rect 14458 27548 14464 27600
rect 14516 27548 14522 27600
rect 14642 27548 14648 27600
rect 14700 27548 14706 27600
rect 15930 27588 15936 27600
rect 15891 27560 15936 27588
rect 15930 27548 15936 27560
rect 15988 27548 15994 27600
rect 16390 27548 16396 27600
rect 16448 27588 16454 27600
rect 16669 27591 16727 27597
rect 16669 27588 16681 27591
rect 16448 27560 16681 27588
rect 16448 27548 16454 27560
rect 16669 27557 16681 27560
rect 16715 27557 16727 27591
rect 16669 27551 16727 27557
rect 12529 27523 12587 27529
rect 11808 27492 12480 27520
rect 4755 27424 5488 27452
rect 4755 27421 4767 27424
rect 4709 27415 4767 27421
rect 5534 27412 5540 27464
rect 5592 27452 5598 27464
rect 5994 27452 6000 27464
rect 5592 27424 6000 27452
rect 5592 27412 5598 27424
rect 5994 27412 6000 27424
rect 6052 27452 6058 27464
rect 6733 27455 6791 27461
rect 6733 27452 6745 27455
rect 6052 27424 6745 27452
rect 6052 27412 6058 27424
rect 6733 27421 6745 27424
rect 6779 27421 6791 27455
rect 6733 27415 6791 27421
rect 7193 27455 7251 27461
rect 7193 27421 7205 27455
rect 7239 27452 7251 27455
rect 8478 27452 8484 27464
rect 7239 27424 8484 27452
rect 7239 27421 7251 27424
rect 7193 27415 7251 27421
rect 8478 27412 8484 27424
rect 8536 27412 8542 27464
rect 9306 27412 9312 27464
rect 9364 27452 9370 27464
rect 10134 27452 10140 27464
rect 9364 27424 10140 27452
rect 9364 27412 9370 27424
rect 10134 27412 10140 27424
rect 10192 27412 10198 27464
rect 10433 27455 10491 27461
rect 10433 27421 10445 27455
rect 10479 27452 10491 27455
rect 10962 27452 10968 27464
rect 10479 27424 10968 27452
rect 10479 27421 10491 27424
rect 10433 27415 10491 27421
rect 10962 27412 10968 27424
rect 11020 27412 11026 27464
rect 12158 27412 12164 27464
rect 12216 27452 12222 27464
rect 12253 27455 12311 27461
rect 12253 27452 12265 27455
rect 12216 27424 12265 27452
rect 12216 27412 12222 27424
rect 12253 27421 12265 27424
rect 12299 27421 12311 27455
rect 12452 27452 12480 27492
rect 12529 27489 12541 27523
rect 12575 27520 12587 27523
rect 13078 27520 13084 27532
rect 12575 27492 13084 27520
rect 12575 27489 12587 27492
rect 12529 27483 12587 27489
rect 13078 27480 13084 27492
rect 13136 27480 13142 27532
rect 13357 27523 13415 27529
rect 13357 27489 13369 27523
rect 13403 27520 13415 27523
rect 13814 27520 13820 27532
rect 13403 27492 13820 27520
rect 13403 27489 13415 27492
rect 13357 27483 13415 27489
rect 13814 27480 13820 27492
rect 13872 27480 13878 27532
rect 14476 27520 14504 27548
rect 14451 27492 14504 27520
rect 14660 27520 14688 27548
rect 15102 27520 15108 27532
rect 14660 27492 15108 27520
rect 12618 27452 12624 27464
rect 12452 27424 12624 27452
rect 12253 27415 12311 27421
rect 12618 27412 12624 27424
rect 12676 27412 12682 27464
rect 13170 27452 13176 27464
rect 13131 27424 13176 27452
rect 13170 27412 13176 27424
rect 13228 27412 13234 27464
rect 13446 27452 13452 27464
rect 13407 27424 13452 27452
rect 13446 27412 13452 27424
rect 13504 27412 13510 27464
rect 3145 27387 3203 27393
rect 3145 27353 3157 27387
rect 3191 27384 3203 27387
rect 3602 27384 3608 27396
rect 3191 27356 3608 27384
rect 3191 27353 3203 27356
rect 3145 27347 3203 27353
rect 3602 27344 3608 27356
rect 3660 27344 3666 27396
rect 3786 27344 3792 27396
rect 3844 27384 3850 27396
rect 3844 27356 6408 27384
rect 3844 27344 3850 27356
rect 2317 27319 2375 27325
rect 2317 27285 2329 27319
rect 2363 27316 2375 27319
rect 4706 27316 4712 27328
rect 2363 27288 4712 27316
rect 2363 27285 2375 27288
rect 2317 27279 2375 27285
rect 4706 27276 4712 27288
rect 4764 27276 4770 27328
rect 6380 27316 6408 27356
rect 6454 27344 6460 27396
rect 6512 27393 6518 27396
rect 6512 27384 6524 27393
rect 6512 27356 6557 27384
rect 6512 27347 6524 27356
rect 6512 27344 6518 27347
rect 6638 27344 6644 27396
rect 6696 27384 6702 27396
rect 7438 27387 7496 27393
rect 7438 27384 7450 27387
rect 6696 27356 7450 27384
rect 6696 27344 6702 27356
rect 7438 27353 7450 27356
rect 7484 27353 7496 27387
rect 7438 27347 7496 27353
rect 7558 27344 7564 27396
rect 7616 27384 7622 27396
rect 11882 27384 11888 27396
rect 7616 27356 8616 27384
rect 7616 27344 7622 27356
rect 8386 27316 8392 27328
rect 6380 27288 8392 27316
rect 8386 27276 8392 27288
rect 8444 27276 8450 27328
rect 8588 27325 8616 27356
rect 9324 27356 11888 27384
rect 8573 27319 8631 27325
rect 8573 27285 8585 27319
rect 8619 27285 8631 27319
rect 8573 27279 8631 27285
rect 8662 27276 8668 27328
rect 8720 27316 8726 27328
rect 9324 27325 9352 27356
rect 11882 27344 11888 27356
rect 11940 27344 11946 27396
rect 12894 27384 12900 27396
rect 11992 27356 12900 27384
rect 9309 27319 9367 27325
rect 9309 27316 9321 27319
rect 8720 27288 9321 27316
rect 8720 27276 8726 27288
rect 9309 27285 9321 27288
rect 9355 27285 9367 27319
rect 9309 27279 9367 27285
rect 9398 27276 9404 27328
rect 9456 27316 9462 27328
rect 11992 27316 12020 27356
rect 12894 27344 12900 27356
rect 12952 27344 12958 27396
rect 13998 27344 14004 27396
rect 14056 27384 14062 27396
rect 14451 27393 14479 27492
rect 15102 27480 15108 27492
rect 15160 27480 15166 27532
rect 15470 27480 15476 27532
rect 15528 27480 15534 27532
rect 15488 27452 15516 27480
rect 14660 27424 15516 27452
rect 14660 27393 14688 27424
rect 15746 27412 15752 27464
rect 15804 27452 15810 27464
rect 16117 27455 16175 27461
rect 16117 27452 16129 27455
rect 15804 27424 16129 27452
rect 15804 27412 15810 27424
rect 16117 27421 16129 27424
rect 16163 27421 16175 27455
rect 16117 27415 16175 27421
rect 16209 27455 16267 27461
rect 16209 27421 16221 27455
rect 16255 27421 16267 27455
rect 16666 27452 16672 27464
rect 16627 27424 16672 27452
rect 16209 27415 16267 27421
rect 14451 27387 14519 27393
rect 14056 27356 14412 27384
rect 14451 27356 14473 27387
rect 14056 27344 14062 27356
rect 9456 27288 12020 27316
rect 9456 27276 9462 27288
rect 12250 27276 12256 27328
rect 12308 27316 12314 27328
rect 12710 27316 12716 27328
rect 12308 27288 12716 27316
rect 12308 27276 12314 27288
rect 12710 27276 12716 27288
rect 12768 27276 12774 27328
rect 12986 27316 12992 27328
rect 12947 27288 12992 27316
rect 12986 27276 12992 27288
rect 13044 27276 13050 27328
rect 13814 27276 13820 27328
rect 13872 27316 13878 27328
rect 14277 27319 14335 27325
rect 14277 27316 14289 27319
rect 13872 27288 14289 27316
rect 13872 27276 13878 27288
rect 14277 27285 14289 27288
rect 14323 27285 14335 27319
rect 14384 27316 14412 27356
rect 14461 27353 14473 27356
rect 14507 27353 14519 27387
rect 14461 27347 14519 27353
rect 14645 27387 14703 27393
rect 14645 27353 14657 27387
rect 14691 27353 14703 27387
rect 15473 27387 15531 27393
rect 14645 27347 14703 27353
rect 15028 27356 15424 27384
rect 15028 27316 15056 27356
rect 14384 27288 15056 27316
rect 14277 27279 14335 27285
rect 15102 27276 15108 27328
rect 15160 27316 15166 27328
rect 15286 27325 15292 27328
rect 15273 27319 15292 27325
rect 15160 27288 15205 27316
rect 15160 27276 15166 27288
rect 15273 27285 15285 27319
rect 15273 27279 15292 27285
rect 15286 27276 15292 27279
rect 15344 27276 15350 27328
rect 15396 27316 15424 27356
rect 15473 27353 15485 27387
rect 15519 27384 15531 27387
rect 15838 27384 15844 27396
rect 15519 27356 15844 27384
rect 15519 27353 15531 27356
rect 15473 27347 15531 27353
rect 15838 27344 15844 27356
rect 15896 27344 15902 27396
rect 15930 27344 15936 27396
rect 15988 27384 15994 27396
rect 16224 27384 16252 27415
rect 16666 27412 16672 27424
rect 16724 27412 16730 27464
rect 16850 27452 16856 27464
rect 16811 27424 16856 27452
rect 16850 27412 16856 27424
rect 16908 27412 16914 27464
rect 28350 27452 28356 27464
rect 28311 27424 28356 27452
rect 28350 27412 28356 27424
rect 28408 27412 28414 27464
rect 17313 27387 17371 27393
rect 17313 27384 17325 27387
rect 15988 27356 16033 27384
rect 16132 27356 17325 27384
rect 15988 27344 15994 27356
rect 16132 27316 16160 27356
rect 17313 27353 17325 27356
rect 17359 27353 17371 27387
rect 17313 27347 17371 27353
rect 15396 27288 16160 27316
rect 1104 27226 29048 27248
rect 1104 27174 7896 27226
rect 7948 27174 7960 27226
rect 8012 27174 8024 27226
rect 8076 27174 8088 27226
rect 8140 27174 8152 27226
rect 8204 27174 14842 27226
rect 14894 27174 14906 27226
rect 14958 27174 14970 27226
rect 15022 27174 15034 27226
rect 15086 27174 15098 27226
rect 15150 27174 21788 27226
rect 21840 27174 21852 27226
rect 21904 27174 21916 27226
rect 21968 27174 21980 27226
rect 22032 27174 22044 27226
rect 22096 27174 28734 27226
rect 28786 27174 28798 27226
rect 28850 27174 28862 27226
rect 28914 27174 28926 27226
rect 28978 27174 28990 27226
rect 29042 27174 29048 27226
rect 1104 27152 29048 27174
rect 1673 27115 1731 27121
rect 1673 27081 1685 27115
rect 1719 27112 1731 27115
rect 2866 27112 2872 27124
rect 1719 27084 2872 27112
rect 1719 27081 1731 27084
rect 1673 27075 1731 27081
rect 2866 27072 2872 27084
rect 2924 27072 2930 27124
rect 3234 27112 3240 27124
rect 3195 27084 3240 27112
rect 3234 27072 3240 27084
rect 3292 27072 3298 27124
rect 3973 27115 4031 27121
rect 3973 27081 3985 27115
rect 4019 27112 4031 27115
rect 6638 27112 6644 27124
rect 4019 27084 6644 27112
rect 4019 27081 4031 27084
rect 3973 27075 4031 27081
rect 6638 27072 6644 27084
rect 6696 27072 6702 27124
rect 8386 27072 8392 27124
rect 8444 27112 8450 27124
rect 10597 27115 10655 27121
rect 10597 27112 10609 27115
rect 8444 27084 10609 27112
rect 8444 27072 8450 27084
rect 10597 27081 10609 27084
rect 10643 27112 10655 27115
rect 10643 27084 12011 27112
rect 10643 27081 10655 27084
rect 10597 27075 10655 27081
rect 5350 27044 5356 27056
rect 1872 27016 5356 27044
rect 1872 26985 1900 27016
rect 5350 27004 5356 27016
rect 5408 27004 5414 27056
rect 5752 27047 5810 27053
rect 5752 27013 5764 27047
rect 5798 27044 5810 27047
rect 7190 27044 7196 27056
rect 5798 27016 7196 27044
rect 5798 27013 5810 27016
rect 5752 27007 5810 27013
rect 7190 27004 7196 27016
rect 7248 27004 7254 27056
rect 8757 27047 8815 27053
rect 8757 27013 8769 27047
rect 8803 27044 8815 27047
rect 9766 27044 9772 27056
rect 8803 27016 9772 27044
rect 8803 27013 8815 27016
rect 8757 27007 8815 27013
rect 9766 27004 9772 27016
rect 9824 27004 9830 27056
rect 10134 27004 10140 27056
rect 10192 27044 10198 27056
rect 11057 27047 11115 27053
rect 11057 27044 11069 27047
rect 10192 27016 11069 27044
rect 10192 27004 10198 27016
rect 11057 27013 11069 27016
rect 11103 27013 11115 27047
rect 11983 27044 12011 27084
rect 12894 27072 12900 27124
rect 12952 27112 12958 27124
rect 12989 27115 13047 27121
rect 12989 27112 13001 27115
rect 12952 27084 13001 27112
rect 12952 27072 12958 27084
rect 12989 27081 13001 27084
rect 13035 27081 13047 27115
rect 12989 27075 13047 27081
rect 13538 27072 13544 27124
rect 13596 27112 13602 27124
rect 13596 27084 14228 27112
rect 13596 27072 13602 27084
rect 13630 27044 13636 27056
rect 11983 27016 13636 27044
rect 11057 27007 11115 27013
rect 1857 26979 1915 26985
rect 1857 26945 1869 26979
rect 1903 26945 1915 26979
rect 1857 26939 1915 26945
rect 2593 26979 2651 26985
rect 2593 26945 2605 26979
rect 2639 26945 2651 26979
rect 2593 26939 2651 26945
rect 1762 26800 1768 26852
rect 1820 26840 1826 26852
rect 2409 26843 2467 26849
rect 2409 26840 2421 26843
rect 1820 26812 2421 26840
rect 1820 26800 1826 26812
rect 2409 26809 2421 26812
rect 2455 26809 2467 26843
rect 2608 26840 2636 26939
rect 2866 26936 2872 26988
rect 2924 26976 2930 26988
rect 3050 26976 3056 26988
rect 2924 26948 3056 26976
rect 2924 26936 2930 26948
rect 3050 26936 3056 26948
rect 3108 26976 3114 26988
rect 3145 26979 3203 26985
rect 3145 26976 3157 26979
rect 3108 26948 3157 26976
rect 3108 26936 3114 26948
rect 3145 26945 3157 26948
rect 3191 26945 3203 26979
rect 3145 26939 3203 26945
rect 3421 26979 3479 26985
rect 3421 26945 3433 26979
rect 3467 26976 3479 26979
rect 3786 26976 3792 26988
rect 3467 26948 3792 26976
rect 3467 26945 3479 26948
rect 3421 26939 3479 26945
rect 3786 26936 3792 26948
rect 3844 26936 3850 26988
rect 3881 26979 3939 26985
rect 3881 26945 3893 26979
rect 3927 26976 3939 26979
rect 3970 26976 3976 26988
rect 3927 26948 3976 26976
rect 3927 26945 3939 26948
rect 3881 26939 3939 26945
rect 3970 26936 3976 26948
rect 4028 26936 4034 26988
rect 4065 26979 4123 26985
rect 4065 26945 4077 26979
rect 4111 26976 4123 26979
rect 4154 26976 4160 26988
rect 4111 26948 4160 26976
rect 4111 26945 4123 26948
rect 4065 26939 4123 26945
rect 4154 26936 4160 26948
rect 4212 26936 4218 26988
rect 5994 26936 6000 26988
rect 6052 26976 6058 26988
rect 6052 26948 6097 26976
rect 6052 26936 6058 26948
rect 6362 26936 6368 26988
rect 6420 26976 6426 26988
rect 7662 26979 7720 26985
rect 7662 26976 7674 26979
rect 6420 26948 7674 26976
rect 6420 26936 6426 26948
rect 7662 26945 7674 26948
rect 7708 26945 7720 26979
rect 7662 26939 7720 26945
rect 7929 26979 7987 26985
rect 7929 26945 7941 26979
rect 7975 26976 7987 26979
rect 8478 26976 8484 26988
rect 7975 26948 8484 26976
rect 7975 26945 7987 26948
rect 7929 26939 7987 26945
rect 8478 26936 8484 26948
rect 8536 26936 8542 26988
rect 8570 26936 8576 26988
rect 8628 26976 8634 26988
rect 8628 26948 8673 26976
rect 8628 26936 8634 26948
rect 8938 26936 8944 26988
rect 8996 26976 9002 26988
rect 9473 26979 9531 26985
rect 9473 26976 9485 26979
rect 8996 26948 9485 26976
rect 8996 26936 9002 26948
rect 9473 26945 9485 26948
rect 9519 26945 9531 26979
rect 9473 26939 9531 26945
rect 6086 26868 6092 26920
rect 6144 26908 6150 26920
rect 8386 26908 8392 26920
rect 6144 26880 6868 26908
rect 8347 26880 8392 26908
rect 6144 26868 6150 26880
rect 2608 26812 4752 26840
rect 2409 26803 2467 26809
rect 3418 26772 3424 26784
rect 3379 26744 3424 26772
rect 3418 26732 3424 26744
rect 3476 26732 3482 26784
rect 4154 26732 4160 26784
rect 4212 26772 4218 26784
rect 4617 26775 4675 26781
rect 4617 26772 4629 26775
rect 4212 26744 4629 26772
rect 4212 26732 4218 26744
rect 4617 26741 4629 26744
rect 4663 26741 4675 26775
rect 4724 26772 4752 26812
rect 5994 26800 6000 26852
rect 6052 26840 6058 26852
rect 6730 26840 6736 26852
rect 6052 26812 6736 26840
rect 6052 26800 6058 26812
rect 6730 26800 6736 26812
rect 6788 26800 6794 26852
rect 6549 26775 6607 26781
rect 6549 26772 6561 26775
rect 4724 26744 6561 26772
rect 4617 26735 4675 26741
rect 6549 26741 6561 26744
rect 6595 26741 6607 26775
rect 6840 26772 6868 26880
rect 8386 26868 8392 26880
rect 8444 26868 8450 26920
rect 8496 26908 8524 26936
rect 9122 26908 9128 26920
rect 8496 26880 9128 26908
rect 9122 26868 9128 26880
rect 9180 26908 9186 26920
rect 9217 26911 9275 26917
rect 9217 26908 9229 26911
rect 9180 26880 9229 26908
rect 9180 26868 9186 26880
rect 9217 26877 9229 26880
rect 9263 26877 9275 26911
rect 9217 26871 9275 26877
rect 10686 26868 10692 26920
rect 10744 26908 10750 26920
rect 10962 26908 10968 26920
rect 10744 26880 10968 26908
rect 10744 26868 10750 26880
rect 10962 26868 10968 26880
rect 11020 26868 11026 26920
rect 11072 26908 11100 27007
rect 13630 27004 13636 27016
rect 13688 27044 13694 27056
rect 13909 27047 13967 27053
rect 13909 27044 13921 27047
rect 13688 27016 13921 27044
rect 13688 27004 13694 27016
rect 13909 27013 13921 27016
rect 13955 27013 13967 27047
rect 13909 27007 13967 27013
rect 13998 27004 14004 27056
rect 14056 27044 14062 27056
rect 14109 27047 14167 27053
rect 14109 27044 14121 27047
rect 14056 27016 14121 27044
rect 14056 27004 14062 27016
rect 14109 27013 14121 27016
rect 14155 27013 14167 27047
rect 14200 27044 14228 27084
rect 14366 27072 14372 27124
rect 14424 27112 14430 27124
rect 14829 27115 14887 27121
rect 14829 27112 14841 27115
rect 14424 27084 14841 27112
rect 14424 27072 14430 27084
rect 14829 27081 14841 27084
rect 14875 27081 14887 27115
rect 14829 27075 14887 27081
rect 15194 27072 15200 27124
rect 15252 27112 15258 27124
rect 15657 27115 15715 27121
rect 15657 27112 15669 27115
rect 15252 27084 15669 27112
rect 15252 27072 15258 27084
rect 15657 27081 15669 27084
rect 15703 27081 15715 27115
rect 15657 27075 15715 27081
rect 15930 27072 15936 27124
rect 15988 27112 15994 27124
rect 16209 27115 16267 27121
rect 16209 27112 16221 27115
rect 15988 27084 16221 27112
rect 15988 27072 15994 27084
rect 16209 27081 16221 27084
rect 16255 27112 16267 27115
rect 17034 27112 17040 27124
rect 16255 27084 17040 27112
rect 16255 27081 16267 27084
rect 16209 27075 16267 27081
rect 17034 27072 17040 27084
rect 17092 27072 17098 27124
rect 14200 27016 15516 27044
rect 14109 27007 14167 27013
rect 11974 26936 11980 26988
rect 12032 26976 12038 26988
rect 13170 26976 13176 26988
rect 12032 26948 12940 26976
rect 13131 26948 13176 26976
rect 12032 26936 12038 26948
rect 12253 26911 12311 26917
rect 11072 26880 11468 26908
rect 9030 26840 9036 26852
rect 7944 26812 9036 26840
rect 7944 26772 7972 26812
rect 9030 26800 9036 26812
rect 9088 26800 9094 26852
rect 6840 26744 7972 26772
rect 6549 26735 6607 26741
rect 8386 26732 8392 26784
rect 8444 26772 8450 26784
rect 10686 26772 10692 26784
rect 8444 26744 10692 26772
rect 8444 26732 8450 26744
rect 10686 26732 10692 26744
rect 10744 26732 10750 26784
rect 11440 26772 11468 26880
rect 12253 26877 12265 26911
rect 12299 26908 12311 26911
rect 12434 26908 12440 26920
rect 12299 26880 12440 26908
rect 12299 26877 12311 26880
rect 12253 26871 12311 26877
rect 12434 26868 12440 26880
rect 12492 26868 12498 26920
rect 12529 26911 12587 26917
rect 12529 26877 12541 26911
rect 12575 26908 12587 26911
rect 12802 26908 12808 26920
rect 12575 26880 12808 26908
rect 12575 26877 12587 26880
rect 12529 26871 12587 26877
rect 12802 26868 12808 26880
rect 12860 26868 12866 26920
rect 12912 26908 12940 26948
rect 13170 26936 13176 26948
rect 13228 26936 13234 26988
rect 13357 26979 13415 26985
rect 13357 26945 13369 26979
rect 13403 26976 13415 26979
rect 14458 26976 14464 26988
rect 13403 26948 14464 26976
rect 13403 26945 13415 26948
rect 13357 26939 13415 26945
rect 14458 26936 14464 26948
rect 14516 26936 14522 26988
rect 14737 26979 14795 26985
rect 14737 26945 14749 26979
rect 14783 26945 14795 26979
rect 14737 26939 14795 26945
rect 13449 26911 13507 26917
rect 13449 26908 13461 26911
rect 12912 26880 13461 26908
rect 13449 26877 13461 26880
rect 13495 26877 13507 26911
rect 14752 26908 14780 26939
rect 14826 26936 14832 26988
rect 14884 26976 14890 26988
rect 15488 26985 15516 27016
rect 15013 26979 15071 26985
rect 15013 26976 15025 26979
rect 14884 26948 15025 26976
rect 14884 26936 14890 26948
rect 15013 26945 15025 26948
rect 15059 26976 15071 26979
rect 15473 26979 15531 26985
rect 15059 26948 15240 26976
rect 15059 26945 15071 26948
rect 15013 26939 15071 26945
rect 13449 26871 13507 26877
rect 14292 26880 14780 26908
rect 14292 26852 14320 26880
rect 14274 26840 14280 26852
rect 14235 26812 14280 26840
rect 14274 26800 14280 26812
rect 14332 26800 14338 26852
rect 14734 26800 14740 26852
rect 14792 26840 14798 26852
rect 15013 26843 15071 26849
rect 15013 26840 15025 26843
rect 14792 26812 15025 26840
rect 14792 26800 14798 26812
rect 15013 26809 15025 26812
rect 15059 26809 15071 26843
rect 15212 26840 15240 26948
rect 15473 26945 15485 26979
rect 15519 26945 15531 26979
rect 15473 26939 15531 26945
rect 15286 26868 15292 26920
rect 15344 26908 15350 26920
rect 16206 26908 16212 26920
rect 15344 26880 16212 26908
rect 15344 26868 15350 26880
rect 16206 26868 16212 26880
rect 16264 26868 16270 26920
rect 15930 26840 15936 26852
rect 15212 26812 15936 26840
rect 15013 26803 15071 26809
rect 15930 26800 15936 26812
rect 15988 26800 15994 26852
rect 12526 26772 12532 26784
rect 11440 26744 12532 26772
rect 12526 26732 12532 26744
rect 12584 26732 12590 26784
rect 14090 26732 14096 26784
rect 14148 26772 14154 26784
rect 14148 26744 14193 26772
rect 14148 26732 14154 26744
rect 1104 26682 28888 26704
rect 1104 26630 4423 26682
rect 4475 26630 4487 26682
rect 4539 26630 4551 26682
rect 4603 26630 4615 26682
rect 4667 26630 4679 26682
rect 4731 26630 11369 26682
rect 11421 26630 11433 26682
rect 11485 26630 11497 26682
rect 11549 26630 11561 26682
rect 11613 26630 11625 26682
rect 11677 26630 18315 26682
rect 18367 26630 18379 26682
rect 18431 26630 18443 26682
rect 18495 26630 18507 26682
rect 18559 26630 18571 26682
rect 18623 26630 25261 26682
rect 25313 26630 25325 26682
rect 25377 26630 25389 26682
rect 25441 26630 25453 26682
rect 25505 26630 25517 26682
rect 25569 26630 28888 26682
rect 1104 26608 28888 26630
rect 2501 26571 2559 26577
rect 2501 26537 2513 26571
rect 2547 26568 2559 26571
rect 4801 26571 4859 26577
rect 2547 26540 4660 26568
rect 2547 26537 2559 26540
rect 2501 26531 2559 26537
rect 3234 26500 3240 26512
rect 3195 26472 3240 26500
rect 3234 26460 3240 26472
rect 3292 26460 3298 26512
rect 4157 26503 4215 26509
rect 4157 26469 4169 26503
rect 4203 26500 4215 26503
rect 4430 26500 4436 26512
rect 4203 26472 4436 26500
rect 4203 26469 4215 26472
rect 4157 26463 4215 26469
rect 4430 26460 4436 26472
rect 4488 26460 4494 26512
rect 2590 26432 2596 26444
rect 2240 26404 2596 26432
rect 1578 26364 1584 26376
rect 1539 26336 1584 26364
rect 1578 26324 1584 26336
rect 1636 26324 1642 26376
rect 2240 26373 2268 26404
rect 2590 26392 2596 26404
rect 2648 26392 2654 26444
rect 4632 26432 4660 26540
rect 4801 26537 4813 26571
rect 4847 26568 4859 26571
rect 4982 26568 4988 26580
rect 4847 26540 4988 26568
rect 4847 26537 4859 26540
rect 4801 26531 4859 26537
rect 4982 26528 4988 26540
rect 5040 26528 5046 26580
rect 5718 26528 5724 26580
rect 5776 26568 5782 26580
rect 5905 26571 5963 26577
rect 5905 26568 5917 26571
rect 5776 26540 5917 26568
rect 5776 26528 5782 26540
rect 5905 26537 5917 26540
rect 5951 26568 5963 26571
rect 6086 26568 6092 26580
rect 5951 26540 6092 26568
rect 5951 26537 5963 26540
rect 5905 26531 5963 26537
rect 6086 26528 6092 26540
rect 6144 26528 6150 26580
rect 6546 26528 6552 26580
rect 6604 26568 6610 26580
rect 7190 26568 7196 26580
rect 6604 26540 7052 26568
rect 7151 26540 7196 26568
rect 6604 26528 6610 26540
rect 5537 26503 5595 26509
rect 5537 26469 5549 26503
rect 5583 26500 5595 26503
rect 5626 26500 5632 26512
rect 5583 26472 5632 26500
rect 5583 26469 5595 26472
rect 5537 26463 5595 26469
rect 5626 26460 5632 26472
rect 5684 26460 5690 26512
rect 6457 26503 6515 26509
rect 6457 26469 6469 26503
rect 6503 26500 6515 26503
rect 6638 26500 6644 26512
rect 6503 26472 6644 26500
rect 6503 26469 6515 26472
rect 6457 26463 6515 26469
rect 6638 26460 6644 26472
rect 6696 26460 6702 26512
rect 2884 26404 4016 26432
rect 4632 26404 5764 26432
rect 2225 26367 2283 26373
rect 2225 26333 2237 26367
rect 2271 26333 2283 26367
rect 2225 26327 2283 26333
rect 2501 26299 2559 26305
rect 2501 26265 2513 26299
rect 2547 26296 2559 26299
rect 2682 26296 2688 26308
rect 2547 26268 2688 26296
rect 2547 26265 2559 26268
rect 2501 26259 2559 26265
rect 2682 26256 2688 26268
rect 2740 26296 2746 26308
rect 2884 26296 2912 26404
rect 3145 26367 3203 26373
rect 3145 26333 3157 26367
rect 3191 26333 3203 26367
rect 3145 26327 3203 26333
rect 2740 26268 2912 26296
rect 2961 26299 3019 26305
rect 2740 26256 2746 26268
rect 2961 26265 2973 26299
rect 3007 26296 3019 26299
rect 3050 26296 3056 26308
rect 3007 26268 3056 26296
rect 3007 26265 3019 26268
rect 2961 26259 3019 26265
rect 3050 26256 3056 26268
rect 3108 26256 3114 26308
rect 3160 26296 3188 26327
rect 3234 26324 3240 26376
rect 3292 26364 3298 26376
rect 3988 26373 4016 26404
rect 3973 26367 4031 26373
rect 3292 26336 3337 26364
rect 3292 26324 3298 26336
rect 3973 26333 3985 26367
rect 4019 26333 4031 26367
rect 3973 26327 4031 26333
rect 4157 26367 4215 26373
rect 4157 26333 4169 26367
rect 4203 26333 4215 26367
rect 4157 26327 4215 26333
rect 3786 26296 3792 26308
rect 3160 26268 3792 26296
rect 3786 26256 3792 26268
rect 3844 26256 3850 26308
rect 2314 26228 2320 26240
rect 2275 26200 2320 26228
rect 2314 26188 2320 26200
rect 2372 26188 2378 26240
rect 3068 26228 3096 26256
rect 3602 26228 3608 26240
rect 3068 26200 3608 26228
rect 3602 26188 3608 26200
rect 3660 26188 3666 26240
rect 4172 26228 4200 26327
rect 4338 26324 4344 26376
rect 4396 26364 4402 26376
rect 5736 26373 5764 26404
rect 6086 26392 6092 26444
rect 6144 26432 6150 26444
rect 6549 26435 6607 26441
rect 6549 26432 6561 26435
rect 6144 26404 6561 26432
rect 6144 26392 6150 26404
rect 6549 26401 6561 26404
rect 6595 26401 6607 26435
rect 7024 26432 7052 26540
rect 7190 26528 7196 26540
rect 7248 26528 7254 26580
rect 7282 26528 7288 26580
rect 7340 26568 7346 26580
rect 7340 26540 8984 26568
rect 7340 26528 7346 26540
rect 8386 26500 8392 26512
rect 8347 26472 8392 26500
rect 8386 26460 8392 26472
rect 8444 26460 8450 26512
rect 8573 26435 8631 26441
rect 8573 26432 8585 26435
rect 7024 26404 8585 26432
rect 6549 26395 6607 26401
rect 8573 26401 8585 26404
rect 8619 26432 8631 26435
rect 8662 26432 8668 26444
rect 8619 26404 8668 26432
rect 8619 26401 8631 26404
rect 8573 26395 8631 26401
rect 8662 26392 8668 26404
rect 8720 26392 8726 26444
rect 8846 26432 8852 26444
rect 8772 26404 8852 26432
rect 4617 26367 4675 26373
rect 4617 26364 4629 26367
rect 4396 26336 4629 26364
rect 4396 26324 4402 26336
rect 4617 26333 4629 26336
rect 4663 26333 4675 26367
rect 4617 26327 4675 26333
rect 5721 26367 5779 26373
rect 5721 26333 5733 26367
rect 5767 26333 5779 26367
rect 5994 26364 6000 26376
rect 5907 26336 6000 26364
rect 5721 26327 5779 26333
rect 5994 26324 6000 26336
rect 6052 26364 6058 26376
rect 6178 26364 6184 26376
rect 6052 26336 6184 26364
rect 6052 26324 6058 26336
rect 6178 26324 6184 26336
rect 6236 26324 6242 26376
rect 6270 26324 6276 26376
rect 6328 26364 6334 26376
rect 6457 26367 6515 26373
rect 6457 26364 6469 26367
rect 6328 26336 6469 26364
rect 6328 26324 6334 26336
rect 6457 26333 6469 26336
rect 6503 26364 6515 26367
rect 7466 26364 7472 26376
rect 6503 26336 7472 26364
rect 6503 26333 6515 26336
rect 6457 26327 6515 26333
rect 7466 26324 7472 26336
rect 7524 26324 7530 26376
rect 7650 26324 7656 26376
rect 7708 26364 7714 26376
rect 7745 26367 7803 26373
rect 7745 26364 7757 26367
rect 7708 26336 7757 26364
rect 7708 26324 7714 26336
rect 7745 26333 7757 26336
rect 7791 26333 7803 26367
rect 7745 26327 7803 26333
rect 8297 26367 8355 26373
rect 8297 26333 8309 26367
rect 8343 26364 8355 26367
rect 8772 26364 8800 26404
rect 8846 26392 8852 26404
rect 8904 26392 8910 26444
rect 8343 26336 8800 26364
rect 8956 26364 8984 26540
rect 9030 26528 9036 26580
rect 9088 26568 9094 26580
rect 9490 26568 9496 26580
rect 9088 26540 9496 26568
rect 9088 26528 9094 26540
rect 9490 26528 9496 26540
rect 9548 26528 9554 26580
rect 10042 26528 10048 26580
rect 10100 26568 10106 26580
rect 10962 26568 10968 26580
rect 10100 26540 10968 26568
rect 10100 26528 10106 26540
rect 10962 26528 10968 26540
rect 11020 26568 11026 26580
rect 12342 26568 12348 26580
rect 11020 26540 12348 26568
rect 11020 26528 11026 26540
rect 12342 26528 12348 26540
rect 12400 26528 12406 26580
rect 12710 26528 12716 26580
rect 12768 26568 12774 26580
rect 12805 26571 12863 26577
rect 12805 26568 12817 26571
rect 12768 26540 12817 26568
rect 12768 26528 12774 26540
rect 12805 26537 12817 26540
rect 12851 26537 12863 26571
rect 12805 26531 12863 26537
rect 12989 26571 13047 26577
rect 12989 26537 13001 26571
rect 13035 26568 13047 26571
rect 13630 26568 13636 26580
rect 13035 26540 13636 26568
rect 13035 26537 13047 26540
rect 12989 26531 13047 26537
rect 13630 26528 13636 26540
rect 13688 26528 13694 26580
rect 14090 26528 14096 26580
rect 14148 26568 14154 26580
rect 18230 26568 18236 26580
rect 14148 26540 18236 26568
rect 14148 26528 14154 26540
rect 18230 26528 18236 26540
rect 18288 26528 18294 26580
rect 10594 26460 10600 26512
rect 10652 26500 10658 26512
rect 13725 26503 13783 26509
rect 13725 26500 13737 26503
rect 10652 26472 13737 26500
rect 10652 26460 10658 26472
rect 13725 26469 13737 26472
rect 13771 26469 13783 26503
rect 13725 26463 13783 26469
rect 13906 26460 13912 26512
rect 13964 26500 13970 26512
rect 15286 26500 15292 26512
rect 13964 26472 15292 26500
rect 13964 26460 13970 26472
rect 15286 26460 15292 26472
rect 15344 26460 15350 26512
rect 9122 26432 9128 26444
rect 9083 26404 9128 26432
rect 9122 26392 9128 26404
rect 9180 26392 9186 26444
rect 10318 26392 10324 26444
rect 10376 26432 10382 26444
rect 10962 26432 10968 26444
rect 10376 26404 10968 26432
rect 10376 26392 10382 26404
rect 10962 26392 10968 26404
rect 11020 26432 11026 26444
rect 11149 26435 11207 26441
rect 11149 26432 11161 26435
rect 11020 26404 11161 26432
rect 11020 26392 11026 26404
rect 11149 26401 11161 26404
rect 11195 26401 11207 26435
rect 11149 26395 11207 26401
rect 11238 26392 11244 26444
rect 11296 26432 11302 26444
rect 11701 26435 11759 26441
rect 11701 26432 11713 26435
rect 11296 26404 11713 26432
rect 11296 26392 11302 26404
rect 11701 26401 11713 26404
rect 11747 26401 11759 26435
rect 12069 26435 12127 26441
rect 11701 26395 11759 26401
rect 11808 26404 12020 26432
rect 11330 26364 11336 26376
rect 8956 26336 11336 26364
rect 8343 26333 8355 26336
rect 8297 26327 8355 26333
rect 11330 26324 11336 26336
rect 11388 26324 11394 26376
rect 6730 26256 6736 26308
rect 6788 26296 6794 26308
rect 8570 26296 8576 26308
rect 6788 26268 6833 26296
rect 8531 26268 8576 26296
rect 6788 26256 6794 26268
rect 8570 26256 8576 26268
rect 8628 26256 8634 26308
rect 8938 26256 8944 26308
rect 8996 26296 9002 26308
rect 9370 26299 9428 26305
rect 9370 26296 9382 26299
rect 8996 26268 9382 26296
rect 8996 26256 9002 26268
rect 9370 26265 9382 26268
rect 9416 26265 9428 26299
rect 11698 26296 11704 26308
rect 9370 26259 9428 26265
rect 9488 26268 11704 26296
rect 6270 26228 6276 26240
rect 4172 26200 6276 26228
rect 6270 26188 6276 26200
rect 6328 26228 6334 26240
rect 7282 26228 7288 26240
rect 6328 26200 7288 26228
rect 6328 26188 6334 26200
rect 7282 26188 7288 26200
rect 7340 26188 7346 26240
rect 9122 26188 9128 26240
rect 9180 26228 9186 26240
rect 9488 26228 9516 26268
rect 11698 26256 11704 26268
rect 11756 26256 11762 26308
rect 9180 26200 9516 26228
rect 9180 26188 9186 26200
rect 9674 26188 9680 26240
rect 9732 26228 9738 26240
rect 10505 26231 10563 26237
rect 10505 26228 10517 26231
rect 9732 26200 10517 26228
rect 9732 26188 9738 26200
rect 10505 26197 10517 26200
rect 10551 26197 10563 26231
rect 10505 26191 10563 26197
rect 10962 26188 10968 26240
rect 11020 26228 11026 26240
rect 11808 26228 11836 26404
rect 11885 26367 11943 26373
rect 11885 26333 11897 26367
rect 11931 26333 11943 26367
rect 11992 26364 12020 26404
rect 12069 26401 12081 26435
rect 12115 26432 12127 26435
rect 12115 26404 12434 26432
rect 12115 26401 12127 26404
rect 12069 26395 12127 26401
rect 12406 26376 12434 26404
rect 12526 26392 12532 26444
rect 12584 26432 12590 26444
rect 13446 26432 13452 26444
rect 12584 26404 13452 26432
rect 12584 26392 12590 26404
rect 13446 26392 13452 26404
rect 13504 26392 13510 26444
rect 13630 26432 13636 26444
rect 13591 26404 13636 26432
rect 13630 26392 13636 26404
rect 13688 26392 13694 26444
rect 16114 26432 16120 26444
rect 13740 26404 16120 26432
rect 12161 26367 12219 26373
rect 12161 26364 12173 26367
rect 11992 26336 12173 26364
rect 11885 26327 11943 26333
rect 12161 26333 12173 26336
rect 12207 26333 12219 26367
rect 12406 26336 12440 26376
rect 12161 26327 12219 26333
rect 11900 26296 11928 26327
rect 12434 26324 12440 26336
rect 12492 26324 12498 26376
rect 13740 26373 13768 26404
rect 16114 26392 16120 26404
rect 16172 26392 16178 26444
rect 13725 26367 13783 26373
rect 12728 26336 13584 26364
rect 11900 26268 12296 26296
rect 11020 26200 11836 26228
rect 12268 26228 12296 26268
rect 12342 26256 12348 26308
rect 12400 26296 12406 26308
rect 12621 26299 12679 26305
rect 12621 26296 12633 26299
rect 12400 26268 12633 26296
rect 12400 26256 12406 26268
rect 12621 26265 12633 26268
rect 12667 26265 12679 26299
rect 12621 26259 12679 26265
rect 12728 26228 12756 26336
rect 12837 26299 12895 26305
rect 12837 26265 12849 26299
rect 12883 26296 12895 26299
rect 13078 26296 13084 26308
rect 12883 26268 13084 26296
rect 12883 26265 12895 26268
rect 12837 26259 12895 26265
rect 13078 26256 13084 26268
rect 13136 26256 13142 26308
rect 13354 26256 13360 26308
rect 13412 26296 13418 26308
rect 13449 26299 13507 26305
rect 13449 26296 13461 26299
rect 13412 26268 13461 26296
rect 13412 26256 13418 26268
rect 13449 26265 13461 26268
rect 13495 26265 13507 26299
rect 13556 26296 13584 26336
rect 13725 26333 13737 26367
rect 13771 26333 13783 26367
rect 13725 26327 13783 26333
rect 14182 26324 14188 26376
rect 14240 26364 14246 26376
rect 14277 26367 14335 26373
rect 14277 26364 14289 26367
rect 14240 26336 14289 26364
rect 14240 26324 14246 26336
rect 14277 26333 14289 26336
rect 14323 26333 14335 26367
rect 14458 26364 14464 26376
rect 14419 26336 14464 26364
rect 14277 26327 14335 26333
rect 14458 26324 14464 26336
rect 14516 26324 14522 26376
rect 17586 26364 17592 26376
rect 14568 26336 17592 26364
rect 14568 26296 14596 26336
rect 17586 26324 17592 26336
rect 17644 26324 17650 26376
rect 14921 26299 14979 26305
rect 14921 26296 14933 26299
rect 13556 26268 14596 26296
rect 14660 26268 14933 26296
rect 13449 26259 13507 26265
rect 12268 26200 12756 26228
rect 11020 26188 11026 26200
rect 13170 26188 13176 26240
rect 13228 26228 13234 26240
rect 14369 26231 14427 26237
rect 14369 26228 14381 26231
rect 13228 26200 14381 26228
rect 13228 26188 13234 26200
rect 14369 26197 14381 26200
rect 14415 26197 14427 26231
rect 14369 26191 14427 26197
rect 14458 26188 14464 26240
rect 14516 26228 14522 26240
rect 14660 26228 14688 26268
rect 14921 26265 14933 26268
rect 14967 26265 14979 26299
rect 14921 26259 14979 26265
rect 15470 26228 15476 26240
rect 14516 26200 14688 26228
rect 15431 26200 15476 26228
rect 14516 26188 14522 26200
rect 15470 26188 15476 26200
rect 15528 26188 15534 26240
rect 1104 26138 29048 26160
rect 1104 26086 7896 26138
rect 7948 26086 7960 26138
rect 8012 26086 8024 26138
rect 8076 26086 8088 26138
rect 8140 26086 8152 26138
rect 8204 26086 14842 26138
rect 14894 26086 14906 26138
rect 14958 26086 14970 26138
rect 15022 26086 15034 26138
rect 15086 26086 15098 26138
rect 15150 26086 21788 26138
rect 21840 26086 21852 26138
rect 21904 26086 21916 26138
rect 21968 26086 21980 26138
rect 22032 26086 22044 26138
rect 22096 26086 28734 26138
rect 28786 26086 28798 26138
rect 28850 26086 28862 26138
rect 28914 26086 28926 26138
rect 28978 26086 28990 26138
rect 29042 26086 29048 26138
rect 1104 26064 29048 26086
rect 1670 26024 1676 26036
rect 1631 25996 1676 26024
rect 1670 25984 1676 25996
rect 1728 25984 1734 26036
rect 4890 25984 4896 26036
rect 4948 26024 4954 26036
rect 7193 26027 7251 26033
rect 4948 25996 6408 26024
rect 4948 25984 4954 25996
rect 4154 25956 4160 25968
rect 1872 25928 4160 25956
rect 1872 25897 1900 25928
rect 4154 25916 4160 25928
rect 4212 25916 4218 25968
rect 5626 25916 5632 25968
rect 5684 25956 5690 25968
rect 5997 25959 6055 25965
rect 5997 25956 6009 25959
rect 5684 25928 6009 25956
rect 5684 25916 5690 25928
rect 5997 25925 6009 25928
rect 6043 25925 6055 25959
rect 6380 25956 6408 25996
rect 7193 25993 7205 26027
rect 7239 25993 7251 26027
rect 7193 25987 7251 25993
rect 8297 26027 8355 26033
rect 8297 25993 8309 26027
rect 8343 26024 8355 26027
rect 8478 26024 8484 26036
rect 8343 25996 8484 26024
rect 8343 25993 8355 25996
rect 8297 25987 8355 25993
rect 6546 25956 6552 25968
rect 6380 25928 6552 25956
rect 5997 25919 6055 25925
rect 6546 25916 6552 25928
rect 6604 25916 6610 25968
rect 1857 25891 1915 25897
rect 1857 25857 1869 25891
rect 1903 25857 1915 25891
rect 1857 25851 1915 25857
rect 3878 25848 3884 25900
rect 3936 25888 3942 25900
rect 3973 25891 4031 25897
rect 3973 25888 3985 25891
rect 3936 25860 3985 25888
rect 3936 25848 3942 25860
rect 3973 25857 3985 25860
rect 4019 25857 4031 25891
rect 3973 25851 4031 25857
rect 5534 25848 5540 25900
rect 5592 25888 5598 25900
rect 5721 25891 5779 25897
rect 5721 25888 5733 25891
rect 5592 25860 5733 25888
rect 5592 25848 5598 25860
rect 5721 25857 5733 25860
rect 5767 25857 5779 25891
rect 5721 25851 5779 25857
rect 5813 25891 5871 25897
rect 5813 25857 5825 25891
rect 5859 25888 5871 25891
rect 6178 25888 6184 25900
rect 5859 25860 6184 25888
rect 5859 25857 5871 25860
rect 5813 25851 5871 25857
rect 6178 25848 6184 25860
rect 6236 25848 6242 25900
rect 6270 25848 6276 25900
rect 6328 25888 6334 25900
rect 7101 25891 7159 25897
rect 7101 25888 7113 25891
rect 6328 25860 7113 25888
rect 6328 25848 6334 25860
rect 7101 25857 7113 25860
rect 7147 25857 7159 25891
rect 7208 25894 7236 25987
rect 8478 25984 8484 25996
rect 8536 25984 8542 26036
rect 10502 26024 10508 26036
rect 10463 25996 10508 26024
rect 10502 25984 10508 25996
rect 10560 25984 10566 26036
rect 10962 26024 10968 26036
rect 10923 25996 10968 26024
rect 10962 25984 10968 25996
rect 11020 25984 11026 26036
rect 11330 25984 11336 26036
rect 11388 26024 11394 26036
rect 12158 26024 12164 26036
rect 11388 25996 12164 26024
rect 11388 25984 11394 25996
rect 12158 25984 12164 25996
rect 12216 26024 12222 26036
rect 12789 26027 12847 26033
rect 12789 26024 12801 26027
rect 12216 25996 12801 26024
rect 12216 25984 12222 25996
rect 12789 25993 12801 25996
rect 12835 26024 12847 26027
rect 12835 25996 14136 26024
rect 12835 25993 12847 25996
rect 12789 25987 12847 25993
rect 9582 25956 9588 25968
rect 9543 25928 9588 25956
rect 9582 25916 9588 25928
rect 9640 25916 9646 25968
rect 11698 25956 11704 25968
rect 11659 25928 11704 25956
rect 11698 25916 11704 25928
rect 11756 25916 11762 25968
rect 12618 25956 12624 25968
rect 11808 25928 12624 25956
rect 7208 25866 7328 25894
rect 7101 25851 7159 25857
rect 14 25780 20 25832
rect 72 25820 78 25832
rect 2961 25823 3019 25829
rect 2961 25820 2973 25823
rect 72 25792 2973 25820
rect 72 25780 78 25792
rect 2961 25789 2973 25792
rect 3007 25789 3019 25823
rect 2961 25783 3019 25789
rect 5077 25823 5135 25829
rect 5077 25789 5089 25823
rect 5123 25820 5135 25823
rect 6914 25820 6920 25832
rect 5123 25792 6920 25820
rect 5123 25789 5135 25792
rect 5077 25783 5135 25789
rect 6914 25780 6920 25792
rect 6972 25780 6978 25832
rect 7006 25780 7012 25832
rect 7064 25820 7070 25832
rect 7300 25820 7328 25866
rect 7377 25891 7435 25897
rect 7377 25857 7389 25891
rect 7423 25888 7435 25891
rect 9858 25888 9864 25900
rect 7423 25860 9864 25888
rect 7423 25857 7435 25860
rect 7377 25851 7435 25857
rect 9858 25848 9864 25860
rect 9916 25848 9922 25900
rect 10042 25888 10048 25900
rect 10003 25860 10048 25888
rect 10042 25848 10048 25860
rect 10100 25848 10106 25900
rect 10318 25888 10324 25900
rect 10279 25860 10324 25888
rect 10318 25848 10324 25860
rect 10376 25848 10382 25900
rect 11808 25888 11836 25928
rect 12618 25916 12624 25928
rect 12676 25916 12682 25968
rect 12986 25956 12992 25968
rect 12947 25928 12992 25956
rect 12986 25916 12992 25928
rect 13044 25916 13050 25968
rect 14108 25956 14136 25996
rect 14734 25956 14740 25968
rect 14108 25928 14228 25956
rect 14695 25928 14740 25956
rect 10428 25860 11836 25888
rect 11885 25891 11943 25897
rect 10428 25820 10456 25860
rect 11885 25857 11897 25891
rect 11931 25888 11943 25891
rect 13170 25888 13176 25900
rect 11931 25860 13176 25888
rect 11931 25857 11943 25860
rect 11885 25851 11943 25857
rect 13170 25848 13176 25860
rect 13228 25848 13234 25900
rect 13437 25891 13495 25897
rect 13437 25888 13449 25891
rect 13372 25860 13449 25888
rect 7064 25792 10456 25820
rect 7064 25780 7070 25792
rect 11146 25780 11152 25832
rect 11204 25820 11210 25832
rect 12161 25823 12219 25829
rect 12161 25820 12173 25823
rect 11204 25792 12173 25820
rect 11204 25780 11210 25792
rect 12161 25789 12173 25792
rect 12207 25789 12219 25823
rect 12161 25783 12219 25789
rect 13078 25780 13084 25832
rect 13136 25820 13142 25832
rect 13372 25820 13400 25860
rect 13437 25857 13449 25860
rect 13483 25857 13495 25891
rect 13437 25851 13495 25857
rect 13538 25848 13544 25900
rect 13596 25888 13602 25900
rect 13633 25891 13691 25897
rect 13633 25888 13645 25891
rect 13596 25860 13645 25888
rect 13596 25848 13602 25860
rect 13633 25857 13645 25860
rect 13679 25888 13691 25891
rect 13906 25888 13912 25900
rect 13679 25860 13912 25888
rect 13679 25857 13691 25860
rect 13633 25851 13691 25857
rect 13906 25848 13912 25860
rect 13964 25848 13970 25900
rect 14200 25888 14228 25928
rect 14734 25916 14740 25928
rect 14792 25916 14798 25968
rect 15378 25888 15384 25900
rect 14200 25860 15384 25888
rect 15378 25848 15384 25860
rect 15436 25848 15442 25900
rect 17126 25888 17132 25900
rect 17087 25860 17132 25888
rect 17126 25848 17132 25860
rect 17184 25888 17190 25900
rect 17589 25891 17647 25897
rect 17589 25888 17601 25891
rect 17184 25860 17601 25888
rect 17184 25848 17190 25860
rect 17589 25857 17601 25860
rect 17635 25857 17647 25891
rect 17589 25851 17647 25857
rect 14093 25823 14151 25829
rect 14093 25820 14105 25823
rect 13136 25792 14105 25820
rect 13136 25780 13142 25792
rect 14093 25789 14105 25792
rect 14139 25820 14151 25823
rect 15470 25820 15476 25832
rect 14139 25792 15476 25820
rect 14139 25789 14151 25792
rect 14093 25783 14151 25789
rect 15470 25780 15476 25792
rect 15528 25820 15534 25832
rect 15528 25792 16988 25820
rect 15528 25780 15534 25792
rect 2130 25712 2136 25764
rect 2188 25752 2194 25764
rect 4982 25752 4988 25764
rect 2188 25724 4988 25752
rect 2188 25712 2194 25724
rect 4982 25712 4988 25724
rect 5040 25712 5046 25764
rect 5997 25755 6055 25761
rect 5997 25721 6009 25755
rect 6043 25752 6055 25755
rect 6086 25752 6092 25764
rect 6043 25724 6092 25752
rect 6043 25721 6055 25724
rect 5997 25715 6055 25721
rect 6086 25712 6092 25724
rect 6144 25712 6150 25764
rect 7190 25712 7196 25764
rect 7248 25752 7254 25764
rect 7377 25755 7435 25761
rect 7377 25752 7389 25755
rect 7248 25724 7389 25752
rect 7248 25712 7254 25724
rect 7377 25721 7389 25724
rect 7423 25721 7435 25755
rect 7377 25715 7435 25721
rect 7834 25712 7840 25764
rect 7892 25752 7898 25764
rect 9306 25752 9312 25764
rect 7892 25724 9312 25752
rect 7892 25712 7898 25724
rect 9306 25712 9312 25724
rect 9364 25712 9370 25764
rect 9858 25712 9864 25764
rect 9916 25752 9922 25764
rect 11054 25752 11060 25764
rect 9916 25724 11060 25752
rect 9916 25712 9922 25724
rect 11054 25712 11060 25724
rect 11112 25712 11118 25764
rect 11974 25752 11980 25764
rect 11900 25724 11980 25752
rect 2314 25684 2320 25696
rect 2275 25656 2320 25684
rect 2314 25644 2320 25656
rect 2372 25644 2378 25696
rect 4062 25644 4068 25696
rect 4120 25684 4126 25696
rect 8110 25684 8116 25696
rect 4120 25656 8116 25684
rect 4120 25644 4126 25656
rect 8110 25644 8116 25656
rect 8168 25644 8174 25696
rect 10137 25687 10195 25693
rect 10137 25653 10149 25687
rect 10183 25684 10195 25687
rect 11900 25684 11928 25724
rect 11974 25712 11980 25724
rect 12032 25712 12038 25764
rect 16850 25752 16856 25764
rect 12406 25724 16856 25752
rect 12066 25684 12072 25696
rect 10183 25656 11928 25684
rect 12027 25656 12072 25684
rect 10183 25653 10195 25656
rect 10137 25647 10195 25653
rect 12066 25644 12072 25656
rect 12124 25684 12130 25696
rect 12406 25684 12434 25724
rect 16850 25712 16856 25724
rect 16908 25712 16914 25764
rect 16960 25761 16988 25792
rect 16945 25755 17003 25761
rect 16945 25721 16957 25755
rect 16991 25721 17003 25755
rect 28350 25752 28356 25764
rect 28311 25724 28356 25752
rect 16945 25715 17003 25721
rect 28350 25712 28356 25724
rect 28408 25712 28414 25764
rect 12618 25684 12624 25696
rect 12124 25656 12434 25684
rect 12579 25656 12624 25684
rect 12124 25644 12130 25656
rect 12618 25644 12624 25656
rect 12676 25644 12682 25696
rect 12710 25644 12716 25696
rect 12768 25684 12774 25696
rect 12805 25687 12863 25693
rect 12805 25684 12817 25687
rect 12768 25656 12817 25684
rect 12768 25644 12774 25656
rect 12805 25653 12817 25656
rect 12851 25684 12863 25687
rect 13262 25684 13268 25696
rect 12851 25656 13268 25684
rect 12851 25653 12863 25656
rect 12805 25647 12863 25653
rect 13262 25644 13268 25656
rect 13320 25644 13326 25696
rect 13633 25687 13691 25693
rect 13633 25653 13645 25687
rect 13679 25684 13691 25687
rect 17402 25684 17408 25696
rect 13679 25656 17408 25684
rect 13679 25653 13691 25656
rect 13633 25647 13691 25653
rect 17402 25644 17408 25656
rect 17460 25644 17466 25696
rect 1104 25594 28888 25616
rect 1104 25542 4423 25594
rect 4475 25542 4487 25594
rect 4539 25542 4551 25594
rect 4603 25542 4615 25594
rect 4667 25542 4679 25594
rect 4731 25542 11369 25594
rect 11421 25542 11433 25594
rect 11485 25542 11497 25594
rect 11549 25542 11561 25594
rect 11613 25542 11625 25594
rect 11677 25542 18315 25594
rect 18367 25542 18379 25594
rect 18431 25542 18443 25594
rect 18495 25542 18507 25594
rect 18559 25542 18571 25594
rect 18623 25542 25261 25594
rect 25313 25542 25325 25594
rect 25377 25542 25389 25594
rect 25441 25542 25453 25594
rect 25505 25542 25517 25594
rect 25569 25542 28888 25594
rect 1104 25520 28888 25542
rect 2225 25483 2283 25489
rect 2225 25449 2237 25483
rect 2271 25480 2283 25483
rect 2958 25480 2964 25492
rect 2271 25452 2964 25480
rect 2271 25449 2283 25452
rect 2225 25443 2283 25449
rect 2958 25440 2964 25452
rect 3016 25440 3022 25492
rect 4982 25440 4988 25492
rect 5040 25480 5046 25492
rect 7377 25483 7435 25489
rect 7377 25480 7389 25483
rect 5040 25452 7389 25480
rect 5040 25440 5046 25452
rect 7377 25449 7389 25452
rect 7423 25449 7435 25483
rect 7377 25443 7435 25449
rect 7466 25440 7472 25492
rect 7524 25480 7530 25492
rect 8205 25483 8263 25489
rect 8205 25480 8217 25483
rect 7524 25452 8217 25480
rect 7524 25440 7530 25452
rect 8205 25449 8217 25452
rect 8251 25449 8263 25483
rect 8205 25443 8263 25449
rect 8573 25483 8631 25489
rect 8573 25449 8585 25483
rect 8619 25480 8631 25483
rect 8938 25480 8944 25492
rect 8619 25452 8944 25480
rect 8619 25449 8631 25452
rect 8573 25443 8631 25449
rect 8938 25440 8944 25452
rect 8996 25440 9002 25492
rect 10137 25483 10195 25489
rect 10137 25449 10149 25483
rect 10183 25480 10195 25483
rect 12066 25480 12072 25492
rect 10183 25452 12072 25480
rect 10183 25449 10195 25452
rect 10137 25443 10195 25449
rect 12066 25440 12072 25452
rect 12124 25440 12130 25492
rect 12526 25440 12532 25492
rect 12584 25480 12590 25492
rect 12713 25483 12771 25489
rect 12713 25480 12725 25483
rect 12584 25452 12725 25480
rect 12584 25440 12590 25452
rect 12713 25449 12725 25452
rect 12759 25449 12771 25483
rect 12713 25443 12771 25449
rect 1581 25415 1639 25421
rect 1581 25381 1593 25415
rect 1627 25412 1639 25415
rect 2774 25412 2780 25424
rect 1627 25384 2780 25412
rect 1627 25381 1639 25384
rect 1581 25375 1639 25381
rect 2774 25372 2780 25384
rect 2832 25372 2838 25424
rect 4893 25415 4951 25421
rect 4893 25381 4905 25415
rect 4939 25412 4951 25415
rect 5442 25412 5448 25424
rect 4939 25384 5448 25412
rect 4939 25381 4951 25384
rect 4893 25375 4951 25381
rect 5442 25372 5448 25384
rect 5500 25372 5506 25424
rect 5902 25372 5908 25424
rect 5960 25412 5966 25424
rect 5997 25415 6055 25421
rect 5997 25412 6009 25415
rect 5960 25384 6009 25412
rect 5960 25372 5966 25384
rect 5997 25381 6009 25384
rect 6043 25381 6055 25415
rect 5997 25375 6055 25381
rect 6917 25415 6975 25421
rect 6917 25381 6929 25415
rect 6963 25412 6975 25415
rect 9030 25412 9036 25424
rect 6963 25384 9036 25412
rect 6963 25381 6975 25384
rect 6917 25375 6975 25381
rect 9030 25372 9036 25384
rect 9088 25372 9094 25424
rect 10962 25412 10968 25424
rect 10796 25384 10968 25412
rect 3418 25304 3424 25356
rect 3476 25344 3482 25356
rect 6825 25347 6883 25353
rect 6825 25344 6837 25347
rect 3476 25316 6837 25344
rect 3476 25304 3482 25316
rect 6825 25313 6837 25316
rect 6871 25313 6883 25347
rect 6825 25307 6883 25313
rect 7098 25304 7104 25356
rect 7156 25344 7162 25356
rect 8110 25344 8116 25356
rect 7156 25316 7696 25344
rect 8071 25316 8116 25344
rect 7156 25304 7162 25316
rect 6178 25276 6184 25288
rect 6139 25248 6184 25276
rect 6178 25236 6184 25248
rect 6236 25236 6242 25288
rect 7668 25285 7696 25316
rect 8110 25304 8116 25316
rect 8168 25344 8174 25356
rect 8168 25316 8616 25344
rect 8168 25304 8174 25316
rect 6917 25279 6975 25285
rect 6917 25245 6929 25279
rect 6963 25276 6975 25279
rect 7653 25279 7711 25285
rect 6963 25248 7604 25276
rect 6963 25245 6975 25248
rect 6917 25239 6975 25245
rect 3050 25168 3056 25220
rect 3108 25208 3114 25220
rect 3421 25211 3479 25217
rect 3421 25208 3433 25211
rect 3108 25180 3433 25208
rect 3108 25168 3114 25180
rect 3421 25177 3433 25180
rect 3467 25208 3479 25211
rect 5537 25211 5595 25217
rect 5537 25208 5549 25211
rect 3467 25180 5549 25208
rect 3467 25177 3479 25180
rect 3421 25171 3479 25177
rect 5537 25177 5549 25180
rect 5583 25208 5595 25211
rect 6454 25208 6460 25220
rect 5583 25180 6460 25208
rect 5583 25177 5595 25180
rect 5537 25171 5595 25177
rect 6454 25168 6460 25180
rect 6512 25208 6518 25220
rect 6641 25211 6699 25217
rect 6641 25208 6653 25211
rect 6512 25180 6653 25208
rect 6512 25168 6518 25180
rect 6641 25177 6653 25180
rect 6687 25208 6699 25211
rect 6730 25208 6736 25220
rect 6687 25180 6736 25208
rect 6687 25177 6699 25180
rect 6641 25171 6699 25177
rect 6730 25168 6736 25180
rect 6788 25168 6794 25220
rect 7377 25211 7435 25217
rect 7377 25177 7389 25211
rect 7423 25208 7435 25211
rect 7466 25208 7472 25220
rect 7423 25180 7472 25208
rect 7423 25177 7435 25180
rect 7377 25171 7435 25177
rect 4246 25140 4252 25152
rect 4207 25112 4252 25140
rect 4246 25100 4252 25112
rect 4304 25140 4310 25152
rect 7392 25140 7420 25171
rect 7466 25168 7472 25180
rect 7524 25168 7530 25220
rect 7576 25208 7604 25248
rect 7653 25245 7665 25279
rect 7699 25245 7711 25279
rect 8386 25276 8392 25288
rect 8347 25248 8392 25276
rect 7653 25239 7711 25245
rect 8386 25236 8392 25248
rect 8444 25236 8450 25288
rect 8588 25276 8616 25316
rect 8846 25304 8852 25356
rect 8904 25344 8910 25356
rect 9766 25344 9772 25356
rect 8904 25316 9772 25344
rect 8904 25304 8910 25316
rect 9766 25304 9772 25316
rect 9824 25304 9830 25356
rect 9674 25276 9680 25288
rect 8588 25248 9680 25276
rect 9674 25236 9680 25248
rect 9732 25236 9738 25288
rect 9858 25276 9864 25288
rect 9819 25248 9864 25276
rect 9858 25236 9864 25248
rect 9916 25236 9922 25288
rect 9950 25236 9956 25288
rect 10008 25276 10014 25288
rect 10796 25285 10824 25384
rect 10962 25372 10968 25384
rect 11020 25372 11026 25424
rect 11974 25372 11980 25424
rect 12032 25412 12038 25424
rect 14274 25412 14280 25424
rect 12032 25384 14280 25412
rect 12032 25372 12038 25384
rect 14274 25372 14280 25384
rect 14332 25372 14338 25424
rect 28350 25412 28356 25424
rect 28311 25384 28356 25412
rect 28350 25372 28356 25384
rect 28408 25372 28414 25424
rect 16574 25344 16580 25356
rect 12544 25316 16580 25344
rect 10781 25279 10839 25285
rect 10008 25248 10053 25276
rect 10008 25236 10014 25248
rect 10781 25245 10793 25279
rect 10827 25245 10839 25279
rect 10781 25239 10839 25245
rect 10965 25279 11023 25285
rect 10965 25245 10977 25279
rect 11011 25276 11023 25279
rect 11054 25276 11060 25288
rect 11011 25248 11060 25276
rect 11011 25245 11023 25248
rect 10965 25239 11023 25245
rect 11054 25236 11060 25248
rect 11112 25236 11118 25288
rect 11146 25236 11152 25288
rect 11204 25276 11210 25288
rect 11701 25279 11759 25285
rect 11701 25276 11713 25279
rect 11204 25248 11713 25276
rect 11204 25236 11210 25248
rect 11701 25245 11713 25248
rect 11747 25245 11759 25279
rect 11701 25239 11759 25245
rect 11790 25236 11796 25288
rect 11848 25276 11854 25288
rect 11885 25279 11943 25285
rect 11885 25276 11897 25279
rect 11848 25248 11897 25276
rect 11848 25236 11854 25248
rect 11885 25245 11897 25248
rect 11931 25245 11943 25279
rect 12544 25276 12572 25316
rect 16574 25304 16580 25316
rect 16632 25304 16638 25356
rect 13078 25276 13084 25288
rect 11885 25239 11943 25245
rect 12084 25248 12572 25276
rect 12636 25248 13084 25276
rect 11974 25208 11980 25220
rect 7576 25180 11980 25208
rect 11974 25168 11980 25180
rect 12032 25168 12038 25220
rect 12084 25152 12112 25248
rect 12342 25168 12348 25220
rect 12400 25208 12406 25220
rect 12636 25217 12664 25248
rect 13078 25236 13084 25248
rect 13136 25276 13142 25288
rect 13265 25279 13323 25285
rect 13265 25276 13277 25279
rect 13136 25248 13277 25276
rect 13136 25236 13142 25248
rect 13265 25245 13277 25248
rect 13311 25245 13323 25279
rect 13265 25239 13323 25245
rect 12621 25211 12679 25217
rect 12621 25208 12633 25211
rect 12400 25180 12633 25208
rect 12400 25168 12406 25180
rect 12621 25177 12633 25180
rect 12667 25177 12679 25211
rect 12621 25171 12679 25177
rect 12710 25168 12716 25220
rect 12768 25208 12774 25220
rect 17678 25208 17684 25220
rect 12768 25180 17684 25208
rect 12768 25168 12774 25180
rect 17678 25168 17684 25180
rect 17736 25168 17742 25220
rect 7558 25140 7564 25152
rect 4304 25112 7420 25140
rect 7519 25112 7564 25140
rect 4304 25100 4310 25112
rect 7558 25100 7564 25112
rect 7616 25140 7622 25152
rect 9122 25140 9128 25152
rect 7616 25112 9128 25140
rect 7616 25100 7622 25112
rect 9122 25100 9128 25112
rect 9180 25100 9186 25152
rect 10594 25140 10600 25152
rect 10555 25112 10600 25140
rect 10594 25100 10600 25112
rect 10652 25100 10658 25152
rect 12066 25140 12072 25152
rect 12027 25112 12072 25140
rect 12066 25100 12072 25112
rect 12124 25100 12130 25152
rect 13998 25100 14004 25152
rect 14056 25140 14062 25152
rect 14274 25140 14280 25152
rect 14056 25112 14280 25140
rect 14056 25100 14062 25112
rect 14274 25100 14280 25112
rect 14332 25100 14338 25152
rect 1104 25050 29048 25072
rect 1104 24998 7896 25050
rect 7948 24998 7960 25050
rect 8012 24998 8024 25050
rect 8076 24998 8088 25050
rect 8140 24998 8152 25050
rect 8204 24998 14842 25050
rect 14894 24998 14906 25050
rect 14958 24998 14970 25050
rect 15022 24998 15034 25050
rect 15086 24998 15098 25050
rect 15150 24998 21788 25050
rect 21840 24998 21852 25050
rect 21904 24998 21916 25050
rect 21968 24998 21980 25050
rect 22032 24998 22044 25050
rect 22096 24998 28734 25050
rect 28786 24998 28798 25050
rect 28850 24998 28862 25050
rect 28914 24998 28926 25050
rect 28978 24998 28990 25050
rect 29042 24998 29048 25050
rect 1104 24976 29048 24998
rect 2133 24939 2191 24945
rect 2133 24905 2145 24939
rect 2179 24936 2191 24939
rect 2222 24936 2228 24948
rect 2179 24908 2228 24936
rect 2179 24905 2191 24908
rect 2133 24899 2191 24905
rect 2222 24896 2228 24908
rect 2280 24896 2286 24948
rect 6178 24896 6184 24948
rect 6236 24936 6242 24948
rect 6236 24908 9720 24936
rect 6236 24896 6242 24908
rect 7098 24868 7104 24880
rect 3160 24840 3464 24868
rect 3160 24800 3188 24840
rect 2746 24772 3188 24800
rect 2746 24744 2774 24772
rect 3234 24760 3240 24812
rect 3292 24800 3298 24812
rect 3329 24803 3387 24809
rect 3329 24800 3341 24803
rect 3292 24772 3341 24800
rect 3292 24760 3298 24772
rect 3329 24769 3341 24772
rect 3375 24769 3387 24803
rect 3436 24800 3464 24840
rect 6840 24840 7104 24868
rect 4246 24800 4252 24812
rect 3436 24772 4252 24800
rect 3329 24763 3387 24769
rect 4246 24760 4252 24772
rect 4304 24760 4310 24812
rect 5074 24760 5080 24812
rect 5132 24800 5138 24812
rect 5169 24803 5227 24809
rect 5169 24800 5181 24803
rect 5132 24772 5181 24800
rect 5132 24760 5138 24772
rect 5169 24769 5181 24772
rect 5215 24769 5227 24803
rect 5169 24763 5227 24769
rect 6733 24803 6791 24809
rect 6733 24769 6745 24803
rect 6779 24800 6791 24803
rect 6840 24800 6868 24840
rect 7098 24828 7104 24840
rect 7156 24828 7162 24880
rect 7558 24828 7564 24880
rect 7616 24868 7622 24880
rect 8202 24868 8208 24880
rect 7616 24840 8208 24868
rect 7616 24828 7622 24840
rect 8202 24828 8208 24840
rect 8260 24828 8266 24880
rect 8294 24828 8300 24880
rect 8352 24868 8358 24880
rect 9582 24868 9588 24880
rect 8352 24840 8524 24868
rect 8352 24828 8358 24840
rect 6779 24772 6868 24800
rect 6779 24769 6791 24772
rect 6733 24763 6791 24769
rect 6914 24760 6920 24812
rect 6972 24800 6978 24812
rect 8496 24809 8524 24840
rect 9355 24837 9413 24843
rect 9543 24840 9588 24868
rect 7469 24803 7527 24809
rect 6972 24772 7017 24800
rect 6972 24760 6978 24772
rect 7469 24769 7481 24803
rect 7515 24769 7527 24803
rect 8389 24803 8447 24809
rect 8389 24800 8401 24803
rect 7469 24763 7527 24769
rect 7576 24772 8401 24800
rect 2682 24732 2688 24744
rect 2595 24704 2688 24732
rect 2682 24692 2688 24704
rect 2740 24704 2774 24744
rect 2740 24692 2746 24704
rect 2866 24692 2872 24744
rect 2924 24732 2930 24744
rect 3881 24735 3939 24741
rect 3881 24732 3893 24735
rect 2924 24704 3893 24732
rect 2924 24692 2930 24704
rect 3881 24701 3893 24704
rect 3927 24701 3939 24735
rect 3881 24695 3939 24701
rect 4525 24735 4583 24741
rect 4525 24701 4537 24735
rect 4571 24732 4583 24735
rect 5997 24735 6055 24741
rect 5997 24732 6009 24735
rect 4571 24704 6009 24732
rect 4571 24701 4583 24704
rect 4525 24695 4583 24701
rect 5997 24701 6009 24704
rect 6043 24732 6055 24735
rect 6454 24732 6460 24744
rect 6043 24704 6460 24732
rect 6043 24701 6055 24704
rect 5997 24695 6055 24701
rect 6454 24692 6460 24704
rect 6512 24692 6518 24744
rect 6822 24692 6828 24744
rect 6880 24732 6886 24744
rect 7484 24732 7512 24763
rect 6880 24704 7512 24732
rect 6880 24692 6886 24704
rect 4798 24624 4804 24676
rect 4856 24664 4862 24676
rect 6733 24667 6791 24673
rect 6733 24664 6745 24667
rect 4856 24636 6745 24664
rect 4856 24624 4862 24636
rect 6733 24633 6745 24636
rect 6779 24633 6791 24667
rect 7576 24664 7604 24772
rect 8389 24769 8401 24772
rect 8435 24769 8447 24803
rect 8389 24763 8447 24769
rect 8481 24803 8539 24809
rect 8481 24769 8493 24803
rect 8527 24769 8539 24803
rect 9355 24803 9367 24837
rect 9401 24803 9413 24837
rect 9582 24828 9588 24840
rect 9640 24828 9646 24880
rect 9692 24868 9720 24908
rect 9766 24896 9772 24948
rect 9824 24936 9830 24948
rect 12342 24936 12348 24948
rect 9824 24908 12348 24936
rect 9824 24896 9830 24908
rect 12342 24896 12348 24908
rect 12400 24896 12406 24948
rect 13814 24868 13820 24880
rect 9692 24840 13820 24868
rect 13814 24828 13820 24840
rect 13872 24828 13878 24880
rect 9355 24797 9413 24803
rect 8481 24763 8539 24769
rect 8202 24692 8208 24744
rect 8260 24732 8266 24744
rect 9370 24732 9398 24797
rect 10410 24760 10416 24812
rect 10468 24800 10474 24812
rect 10597 24803 10655 24809
rect 10597 24800 10609 24803
rect 10468 24772 10609 24800
rect 10468 24760 10474 24772
rect 10597 24769 10609 24772
rect 10643 24769 10655 24803
rect 10597 24763 10655 24769
rect 10686 24760 10692 24812
rect 10744 24800 10750 24812
rect 11701 24803 11759 24809
rect 11701 24800 11713 24803
rect 10744 24772 11713 24800
rect 10744 24760 10750 24772
rect 11701 24769 11713 24772
rect 11747 24769 11759 24803
rect 11882 24800 11888 24812
rect 11843 24772 11888 24800
rect 11701 24763 11759 24769
rect 11882 24760 11888 24772
rect 11940 24760 11946 24812
rect 11974 24760 11980 24812
rect 12032 24800 12038 24812
rect 12529 24803 12587 24809
rect 12529 24800 12541 24803
rect 12032 24772 12077 24800
rect 12406 24772 12541 24800
rect 12032 24760 12038 24772
rect 8260 24704 9398 24732
rect 8260 24692 8266 24704
rect 9582 24692 9588 24744
rect 9640 24732 9646 24744
rect 10873 24735 10931 24741
rect 10873 24732 10885 24735
rect 9640 24704 10885 24732
rect 9640 24692 9646 24704
rect 10873 24701 10885 24704
rect 10919 24732 10931 24735
rect 10919 24704 11100 24732
rect 10919 24701 10931 24704
rect 10873 24695 10931 24701
rect 6733 24627 6791 24633
rect 6840 24636 7604 24664
rect 7653 24667 7711 24673
rect 6270 24556 6276 24608
rect 6328 24596 6334 24608
rect 6840 24596 6868 24636
rect 7653 24633 7665 24667
rect 7699 24664 7711 24667
rect 7742 24664 7748 24676
rect 7699 24636 7748 24664
rect 7699 24633 7711 24636
rect 7653 24627 7711 24633
rect 7742 24624 7748 24636
rect 7800 24624 7806 24676
rect 10045 24667 10103 24673
rect 10045 24664 10057 24667
rect 8404 24636 10057 24664
rect 6328 24568 6868 24596
rect 6328 24556 6334 24568
rect 7558 24556 7564 24608
rect 7616 24596 7622 24608
rect 8404 24596 8432 24636
rect 10045 24633 10057 24636
rect 10091 24664 10103 24667
rect 10689 24667 10747 24673
rect 10689 24664 10701 24667
rect 10091 24636 10701 24664
rect 10091 24633 10103 24636
rect 10045 24627 10103 24633
rect 10689 24633 10701 24636
rect 10735 24664 10747 24667
rect 10962 24664 10968 24676
rect 10735 24636 10968 24664
rect 10735 24633 10747 24636
rect 10689 24627 10747 24633
rect 10962 24624 10968 24636
rect 11020 24624 11026 24676
rect 7616 24568 8432 24596
rect 7616 24556 7622 24568
rect 8478 24556 8484 24608
rect 8536 24596 8542 24608
rect 9217 24599 9275 24605
rect 9217 24596 9229 24599
rect 8536 24568 9229 24596
rect 8536 24556 8542 24568
rect 9217 24565 9229 24568
rect 9263 24565 9275 24599
rect 9217 24559 9275 24565
rect 9401 24599 9459 24605
rect 9401 24565 9413 24599
rect 9447 24596 9459 24599
rect 9490 24596 9496 24608
rect 9447 24568 9496 24596
rect 9447 24565 9459 24568
rect 9401 24559 9459 24565
rect 9490 24556 9496 24568
rect 9548 24556 9554 24608
rect 10778 24556 10784 24608
rect 10836 24596 10842 24608
rect 11072 24596 11100 24704
rect 11146 24692 11152 24744
rect 11204 24732 11210 24744
rect 12406 24732 12434 24772
rect 12529 24769 12541 24772
rect 12575 24800 12587 24803
rect 12894 24800 12900 24812
rect 12575 24772 12900 24800
rect 12575 24769 12587 24772
rect 12529 24763 12587 24769
rect 12894 24760 12900 24772
rect 12952 24760 12958 24812
rect 13354 24800 13360 24812
rect 13267 24772 13360 24800
rect 13354 24760 13360 24772
rect 13412 24800 13418 24812
rect 13906 24800 13912 24812
rect 13412 24772 13912 24800
rect 13412 24760 13418 24772
rect 13906 24760 13912 24772
rect 13964 24800 13970 24812
rect 14734 24800 14740 24812
rect 13964 24772 14740 24800
rect 13964 24760 13970 24772
rect 14734 24760 14740 24772
rect 14792 24760 14798 24812
rect 11204 24704 12434 24732
rect 11204 24692 11210 24704
rect 11698 24664 11704 24676
rect 11659 24636 11704 24664
rect 11698 24624 11704 24636
rect 11756 24624 11762 24676
rect 12250 24596 12256 24608
rect 10836 24568 10881 24596
rect 11072 24568 12256 24596
rect 10836 24556 10842 24568
rect 12250 24556 12256 24568
rect 12308 24556 12314 24608
rect 1104 24506 28888 24528
rect 1104 24454 4423 24506
rect 4475 24454 4487 24506
rect 4539 24454 4551 24506
rect 4603 24454 4615 24506
rect 4667 24454 4679 24506
rect 4731 24454 11369 24506
rect 11421 24454 11433 24506
rect 11485 24454 11497 24506
rect 11549 24454 11561 24506
rect 11613 24454 11625 24506
rect 11677 24454 18315 24506
rect 18367 24454 18379 24506
rect 18431 24454 18443 24506
rect 18495 24454 18507 24506
rect 18559 24454 18571 24506
rect 18623 24454 25261 24506
rect 25313 24454 25325 24506
rect 25377 24454 25389 24506
rect 25441 24454 25453 24506
rect 25505 24454 25517 24506
rect 25569 24454 28888 24506
rect 1104 24432 28888 24454
rect 2501 24395 2559 24401
rect 2501 24361 2513 24395
rect 2547 24392 2559 24395
rect 2866 24392 2872 24404
rect 2547 24364 2872 24392
rect 2547 24361 2559 24364
rect 2501 24355 2559 24361
rect 2866 24352 2872 24364
rect 2924 24352 2930 24404
rect 4341 24395 4399 24401
rect 4341 24361 4353 24395
rect 4387 24392 4399 24395
rect 4890 24392 4896 24404
rect 4387 24364 4896 24392
rect 4387 24361 4399 24364
rect 4341 24355 4399 24361
rect 4890 24352 4896 24364
rect 4948 24352 4954 24404
rect 8386 24392 8392 24404
rect 8347 24364 8392 24392
rect 8386 24352 8392 24364
rect 8444 24352 8450 24404
rect 8662 24352 8668 24404
rect 8720 24392 8726 24404
rect 9766 24392 9772 24404
rect 8720 24364 9772 24392
rect 8720 24352 8726 24364
rect 9766 24352 9772 24364
rect 9824 24352 9830 24404
rect 9950 24392 9956 24404
rect 9911 24364 9956 24392
rect 9950 24352 9956 24364
rect 10008 24352 10014 24404
rect 10781 24395 10839 24401
rect 10781 24361 10793 24395
rect 10827 24392 10839 24395
rect 10870 24392 10876 24404
rect 10827 24364 10876 24392
rect 10827 24361 10839 24364
rect 10781 24355 10839 24361
rect 10870 24352 10876 24364
rect 10928 24352 10934 24404
rect 10962 24352 10968 24404
rect 11020 24392 11026 24404
rect 11790 24392 11796 24404
rect 11020 24364 11796 24392
rect 11020 24352 11026 24364
rect 11790 24352 11796 24364
rect 11848 24392 11854 24404
rect 12161 24395 12219 24401
rect 12161 24392 12173 24395
rect 11848 24364 12173 24392
rect 11848 24352 11854 24364
rect 12161 24361 12173 24364
rect 12207 24361 12219 24395
rect 12161 24355 12219 24361
rect 3970 24284 3976 24336
rect 4028 24324 4034 24336
rect 9125 24327 9183 24333
rect 9125 24324 9137 24327
rect 4028 24296 9137 24324
rect 4028 24284 4034 24296
rect 9125 24293 9137 24296
rect 9171 24293 9183 24327
rect 9125 24287 9183 24293
rect 10045 24327 10103 24333
rect 10045 24293 10057 24327
rect 10091 24324 10103 24327
rect 16666 24324 16672 24336
rect 10091 24296 16672 24324
rect 10091 24293 10103 24296
rect 10045 24287 10103 24293
rect 16666 24284 16672 24296
rect 16724 24284 16730 24336
rect 5442 24216 5448 24268
rect 5500 24256 5506 24268
rect 6914 24256 6920 24268
rect 5500 24228 6920 24256
rect 5500 24216 5506 24228
rect 6914 24216 6920 24228
rect 6972 24256 6978 24268
rect 7009 24259 7067 24265
rect 7009 24256 7021 24259
rect 6972 24228 7021 24256
rect 6972 24216 6978 24228
rect 7009 24225 7021 24228
rect 7055 24225 7067 24259
rect 7009 24219 7067 24225
rect 7098 24216 7104 24268
rect 7156 24256 7162 24268
rect 7156 24228 9444 24256
rect 7156 24216 7162 24228
rect 1578 24188 1584 24200
rect 1539 24160 1584 24188
rect 1578 24148 1584 24160
rect 1636 24148 1642 24200
rect 6362 24148 6368 24200
rect 6420 24188 6426 24200
rect 8389 24191 8447 24197
rect 8389 24188 8401 24191
rect 6420 24160 8401 24188
rect 6420 24148 6426 24160
rect 8389 24157 8401 24160
rect 8435 24188 8447 24191
rect 8478 24188 8484 24200
rect 8435 24160 8484 24188
rect 8435 24157 8447 24160
rect 8389 24151 8447 24157
rect 8478 24148 8484 24160
rect 8536 24148 8542 24200
rect 8573 24191 8631 24197
rect 8573 24157 8585 24191
rect 8619 24188 8631 24191
rect 8662 24188 8668 24200
rect 8619 24160 8668 24188
rect 8619 24157 8631 24160
rect 8573 24151 8631 24157
rect 8662 24148 8668 24160
rect 8720 24148 8726 24200
rect 9214 24148 9220 24200
rect 9272 24188 9278 24200
rect 9416 24197 9444 24228
rect 9582 24216 9588 24268
rect 9640 24256 9646 24268
rect 10137 24259 10195 24265
rect 10137 24256 10149 24259
rect 9640 24228 10149 24256
rect 9640 24216 9646 24228
rect 10137 24225 10149 24228
rect 10183 24225 10195 24259
rect 12066 24256 12072 24268
rect 10137 24219 10195 24225
rect 10612 24228 12072 24256
rect 9309 24191 9367 24197
rect 9309 24188 9321 24191
rect 9272 24160 9321 24188
rect 9272 24148 9278 24160
rect 9309 24157 9321 24160
rect 9355 24157 9367 24191
rect 9309 24151 9367 24157
rect 9401 24191 9459 24197
rect 9401 24157 9413 24191
rect 9447 24157 9459 24191
rect 9858 24188 9864 24200
rect 9819 24160 9864 24188
rect 9401 24151 9459 24157
rect 9858 24148 9864 24160
rect 9916 24148 9922 24200
rect 10612 24197 10640 24228
rect 12066 24216 12072 24228
rect 12124 24216 12130 24268
rect 10597 24191 10655 24197
rect 10597 24157 10609 24191
rect 10643 24157 10655 24191
rect 10778 24188 10784 24200
rect 10739 24160 10784 24188
rect 10597 24151 10655 24157
rect 10778 24148 10784 24160
rect 10836 24148 10842 24200
rect 28350 24188 28356 24200
rect 28311 24160 28356 24188
rect 28350 24148 28356 24160
rect 28408 24148 28414 24200
rect 5077 24123 5135 24129
rect 5077 24089 5089 24123
rect 5123 24120 5135 24123
rect 7558 24120 7564 24132
rect 5123 24092 7564 24120
rect 5123 24089 5135 24092
rect 5077 24083 5135 24089
rect 7558 24080 7564 24092
rect 7616 24080 7622 24132
rect 7650 24080 7656 24132
rect 7708 24120 7714 24132
rect 9125 24123 9183 24129
rect 9125 24120 9137 24123
rect 7708 24092 9137 24120
rect 7708 24080 7714 24092
rect 9125 24089 9137 24092
rect 9171 24089 9183 24123
rect 9125 24083 9183 24089
rect 10410 24080 10416 24132
rect 10468 24120 10474 24132
rect 11146 24120 11152 24132
rect 10468 24092 11152 24120
rect 10468 24080 10474 24092
rect 11146 24080 11152 24092
rect 11204 24120 11210 24132
rect 11241 24123 11299 24129
rect 11241 24120 11253 24123
rect 11204 24092 11253 24120
rect 11204 24080 11210 24092
rect 11241 24089 11253 24092
rect 11287 24089 11299 24123
rect 11241 24083 11299 24089
rect 6454 24052 6460 24064
rect 6415 24024 6460 24052
rect 6454 24012 6460 24024
rect 6512 24012 6518 24064
rect 7466 24012 7472 24064
rect 7524 24052 7530 24064
rect 7745 24055 7803 24061
rect 7745 24052 7757 24055
rect 7524 24024 7757 24052
rect 7524 24012 7530 24024
rect 7745 24021 7757 24024
rect 7791 24021 7803 24055
rect 7745 24015 7803 24021
rect 1104 23962 29048 23984
rect 1104 23910 7896 23962
rect 7948 23910 7960 23962
rect 8012 23910 8024 23962
rect 8076 23910 8088 23962
rect 8140 23910 8152 23962
rect 8204 23910 14842 23962
rect 14894 23910 14906 23962
rect 14958 23910 14970 23962
rect 15022 23910 15034 23962
rect 15086 23910 15098 23962
rect 15150 23910 21788 23962
rect 21840 23910 21852 23962
rect 21904 23910 21916 23962
rect 21968 23910 21980 23962
rect 22032 23910 22044 23962
rect 22096 23910 28734 23962
rect 28786 23910 28798 23962
rect 28850 23910 28862 23962
rect 28914 23910 28926 23962
rect 28978 23910 28990 23962
rect 29042 23910 29048 23962
rect 1104 23888 29048 23910
rect 4341 23851 4399 23857
rect 4341 23817 4353 23851
rect 4387 23848 4399 23851
rect 5442 23848 5448 23860
rect 4387 23820 5448 23848
rect 4387 23817 4399 23820
rect 4341 23811 4399 23817
rect 5442 23808 5448 23820
rect 5500 23808 5506 23860
rect 6914 23848 6920 23860
rect 6875 23820 6920 23848
rect 6914 23808 6920 23820
rect 6972 23808 6978 23860
rect 7374 23808 7380 23860
rect 7432 23848 7438 23860
rect 9861 23851 9919 23857
rect 9861 23848 9873 23851
rect 7432 23820 9873 23848
rect 7432 23808 7438 23820
rect 9861 23817 9873 23820
rect 9907 23817 9919 23851
rect 9861 23811 9919 23817
rect 10505 23851 10563 23857
rect 10505 23817 10517 23851
rect 10551 23848 10563 23851
rect 14274 23848 14280 23860
rect 10551 23820 14280 23848
rect 10551 23817 10563 23820
rect 10505 23811 10563 23817
rect 5074 23740 5080 23792
rect 5132 23780 5138 23792
rect 10410 23780 10416 23792
rect 5132 23752 10416 23780
rect 5132 23740 5138 23752
rect 10410 23740 10416 23752
rect 10468 23740 10474 23792
rect 8570 23672 8576 23724
rect 8628 23712 8634 23724
rect 9769 23715 9827 23721
rect 9769 23712 9781 23715
rect 8628 23684 9781 23712
rect 8628 23672 8634 23684
rect 9769 23681 9781 23684
rect 9815 23681 9827 23715
rect 9769 23675 9827 23681
rect 9953 23715 10011 23721
rect 9953 23681 9965 23715
rect 9999 23712 10011 23715
rect 10520 23712 10548 23811
rect 14274 23808 14280 23820
rect 14332 23808 14338 23860
rect 9999 23684 10548 23712
rect 9999 23681 10011 23684
rect 9953 23675 10011 23681
rect 6914 23604 6920 23656
rect 6972 23644 6978 23656
rect 8662 23644 8668 23656
rect 6972 23616 8668 23644
rect 6972 23604 6978 23616
rect 8662 23604 8668 23616
rect 8720 23604 8726 23656
rect 9309 23647 9367 23653
rect 9309 23613 9321 23647
rect 9355 23644 9367 23647
rect 9582 23644 9588 23656
rect 9355 23616 9588 23644
rect 9355 23613 9367 23616
rect 9309 23607 9367 23613
rect 9582 23604 9588 23616
rect 9640 23644 9646 23656
rect 10965 23647 11023 23653
rect 10965 23644 10977 23647
rect 9640 23616 10977 23644
rect 9640 23604 9646 23616
rect 10965 23613 10977 23616
rect 11011 23613 11023 23647
rect 10965 23607 11023 23613
rect 1578 23508 1584 23520
rect 1539 23480 1584 23508
rect 1578 23468 1584 23480
rect 1636 23468 1642 23520
rect 6454 23468 6460 23520
rect 6512 23508 6518 23520
rect 13906 23508 13912 23520
rect 6512 23480 13912 23508
rect 6512 23468 6518 23480
rect 13906 23468 13912 23480
rect 13964 23468 13970 23520
rect 1104 23418 28888 23440
rect 1104 23366 4423 23418
rect 4475 23366 4487 23418
rect 4539 23366 4551 23418
rect 4603 23366 4615 23418
rect 4667 23366 4679 23418
rect 4731 23366 11369 23418
rect 11421 23366 11433 23418
rect 11485 23366 11497 23418
rect 11549 23366 11561 23418
rect 11613 23366 11625 23418
rect 11677 23366 18315 23418
rect 18367 23366 18379 23418
rect 18431 23366 18443 23418
rect 18495 23366 18507 23418
rect 18559 23366 18571 23418
rect 18623 23366 25261 23418
rect 25313 23366 25325 23418
rect 25377 23366 25389 23418
rect 25441 23366 25453 23418
rect 25505 23366 25517 23418
rect 25569 23366 28888 23418
rect 1104 23344 28888 23366
rect 9214 23264 9220 23316
rect 9272 23304 9278 23316
rect 9493 23307 9551 23313
rect 9493 23304 9505 23307
rect 9272 23276 9505 23304
rect 9272 23264 9278 23276
rect 9493 23273 9505 23276
rect 9539 23273 9551 23307
rect 9493 23267 9551 23273
rect 28350 23100 28356 23112
rect 28311 23072 28356 23100
rect 28350 23060 28356 23072
rect 28408 23060 28414 23112
rect 1104 22874 29048 22896
rect 1104 22822 7896 22874
rect 7948 22822 7960 22874
rect 8012 22822 8024 22874
rect 8076 22822 8088 22874
rect 8140 22822 8152 22874
rect 8204 22822 14842 22874
rect 14894 22822 14906 22874
rect 14958 22822 14970 22874
rect 15022 22822 15034 22874
rect 15086 22822 15098 22874
rect 15150 22822 21788 22874
rect 21840 22822 21852 22874
rect 21904 22822 21916 22874
rect 21968 22822 21980 22874
rect 22032 22822 22044 22874
rect 22096 22822 28734 22874
rect 28786 22822 28798 22874
rect 28850 22822 28862 22874
rect 28914 22822 28926 22874
rect 28978 22822 28990 22874
rect 29042 22822 29048 22874
rect 1104 22800 29048 22822
rect 1578 22420 1584 22432
rect 1539 22392 1584 22420
rect 1578 22380 1584 22392
rect 1636 22380 1642 22432
rect 1104 22330 28888 22352
rect 1104 22278 4423 22330
rect 4475 22278 4487 22330
rect 4539 22278 4551 22330
rect 4603 22278 4615 22330
rect 4667 22278 4679 22330
rect 4731 22278 11369 22330
rect 11421 22278 11433 22330
rect 11485 22278 11497 22330
rect 11549 22278 11561 22330
rect 11613 22278 11625 22330
rect 11677 22278 18315 22330
rect 18367 22278 18379 22330
rect 18431 22278 18443 22330
rect 18495 22278 18507 22330
rect 18559 22278 18571 22330
rect 18623 22278 25261 22330
rect 25313 22278 25325 22330
rect 25377 22278 25389 22330
rect 25441 22278 25453 22330
rect 25505 22278 25517 22330
rect 25569 22278 28888 22330
rect 1104 22256 28888 22278
rect 28350 22012 28356 22024
rect 28311 21984 28356 22012
rect 28350 21972 28356 21984
rect 28408 21972 28414 22024
rect 1104 21786 29048 21808
rect 1104 21734 7896 21786
rect 7948 21734 7960 21786
rect 8012 21734 8024 21786
rect 8076 21734 8088 21786
rect 8140 21734 8152 21786
rect 8204 21734 14842 21786
rect 14894 21734 14906 21786
rect 14958 21734 14970 21786
rect 15022 21734 15034 21786
rect 15086 21734 15098 21786
rect 15150 21734 21788 21786
rect 21840 21734 21852 21786
rect 21904 21734 21916 21786
rect 21968 21734 21980 21786
rect 22032 21734 22044 21786
rect 22096 21734 28734 21786
rect 28786 21734 28798 21786
rect 28850 21734 28862 21786
rect 28914 21734 28926 21786
rect 28978 21734 28990 21786
rect 29042 21734 29048 21786
rect 1104 21712 29048 21734
rect 1578 21468 1584 21480
rect 1539 21440 1584 21468
rect 1578 21428 1584 21440
rect 1636 21428 1642 21480
rect 28350 21332 28356 21344
rect 28311 21304 28356 21332
rect 28350 21292 28356 21304
rect 28408 21292 28414 21344
rect 1104 21242 28888 21264
rect 1104 21190 4423 21242
rect 4475 21190 4487 21242
rect 4539 21190 4551 21242
rect 4603 21190 4615 21242
rect 4667 21190 4679 21242
rect 4731 21190 11369 21242
rect 11421 21190 11433 21242
rect 11485 21190 11497 21242
rect 11549 21190 11561 21242
rect 11613 21190 11625 21242
rect 11677 21190 18315 21242
rect 18367 21190 18379 21242
rect 18431 21190 18443 21242
rect 18495 21190 18507 21242
rect 18559 21190 18571 21242
rect 18623 21190 25261 21242
rect 25313 21190 25325 21242
rect 25377 21190 25389 21242
rect 25441 21190 25453 21242
rect 25505 21190 25517 21242
rect 25569 21190 28888 21242
rect 1104 21168 28888 21190
rect 1104 20698 29048 20720
rect 1104 20646 7896 20698
rect 7948 20646 7960 20698
rect 8012 20646 8024 20698
rect 8076 20646 8088 20698
rect 8140 20646 8152 20698
rect 8204 20646 14842 20698
rect 14894 20646 14906 20698
rect 14958 20646 14970 20698
rect 15022 20646 15034 20698
rect 15086 20646 15098 20698
rect 15150 20646 21788 20698
rect 21840 20646 21852 20698
rect 21904 20646 21916 20698
rect 21968 20646 21980 20698
rect 22032 20646 22044 20698
rect 22096 20646 28734 20698
rect 28786 20646 28798 20698
rect 28850 20646 28862 20698
rect 28914 20646 28926 20698
rect 28978 20646 28990 20698
rect 29042 20646 29048 20698
rect 1104 20624 29048 20646
rect 1578 20244 1584 20256
rect 1539 20216 1584 20244
rect 1578 20204 1584 20216
rect 1636 20204 1642 20256
rect 1104 20154 28888 20176
rect 1104 20102 4423 20154
rect 4475 20102 4487 20154
rect 4539 20102 4551 20154
rect 4603 20102 4615 20154
rect 4667 20102 4679 20154
rect 4731 20102 11369 20154
rect 11421 20102 11433 20154
rect 11485 20102 11497 20154
rect 11549 20102 11561 20154
rect 11613 20102 11625 20154
rect 11677 20102 18315 20154
rect 18367 20102 18379 20154
rect 18431 20102 18443 20154
rect 18495 20102 18507 20154
rect 18559 20102 18571 20154
rect 18623 20102 25261 20154
rect 25313 20102 25325 20154
rect 25377 20102 25389 20154
rect 25441 20102 25453 20154
rect 25505 20102 25517 20154
rect 25569 20102 28888 20154
rect 1104 20080 28888 20102
rect 28350 19972 28356 19984
rect 28311 19944 28356 19972
rect 28350 19932 28356 19944
rect 28408 19932 28414 19984
rect 1578 19836 1584 19848
rect 1539 19808 1584 19836
rect 1578 19796 1584 19808
rect 1636 19796 1642 19848
rect 1104 19610 29048 19632
rect 1104 19558 7896 19610
rect 7948 19558 7960 19610
rect 8012 19558 8024 19610
rect 8076 19558 8088 19610
rect 8140 19558 8152 19610
rect 8204 19558 14842 19610
rect 14894 19558 14906 19610
rect 14958 19558 14970 19610
rect 15022 19558 15034 19610
rect 15086 19558 15098 19610
rect 15150 19558 21788 19610
rect 21840 19558 21852 19610
rect 21904 19558 21916 19610
rect 21968 19558 21980 19610
rect 22032 19558 22044 19610
rect 22096 19558 28734 19610
rect 28786 19558 28798 19610
rect 28850 19558 28862 19610
rect 28914 19558 28926 19610
rect 28978 19558 28990 19610
rect 29042 19558 29048 19610
rect 1104 19536 29048 19558
rect 28350 19156 28356 19168
rect 28311 19128 28356 19156
rect 28350 19116 28356 19128
rect 28408 19116 28414 19168
rect 1104 19066 28888 19088
rect 1104 19014 4423 19066
rect 4475 19014 4487 19066
rect 4539 19014 4551 19066
rect 4603 19014 4615 19066
rect 4667 19014 4679 19066
rect 4731 19014 11369 19066
rect 11421 19014 11433 19066
rect 11485 19014 11497 19066
rect 11549 19014 11561 19066
rect 11613 19014 11625 19066
rect 11677 19014 18315 19066
rect 18367 19014 18379 19066
rect 18431 19014 18443 19066
rect 18495 19014 18507 19066
rect 18559 19014 18571 19066
rect 18623 19014 25261 19066
rect 25313 19014 25325 19066
rect 25377 19014 25389 19066
rect 25441 19014 25453 19066
rect 25505 19014 25517 19066
rect 25569 19014 28888 19066
rect 1104 18992 28888 19014
rect 1104 18522 29048 18544
rect 1104 18470 7896 18522
rect 7948 18470 7960 18522
rect 8012 18470 8024 18522
rect 8076 18470 8088 18522
rect 8140 18470 8152 18522
rect 8204 18470 14842 18522
rect 14894 18470 14906 18522
rect 14958 18470 14970 18522
rect 15022 18470 15034 18522
rect 15086 18470 15098 18522
rect 15150 18470 21788 18522
rect 21840 18470 21852 18522
rect 21904 18470 21916 18522
rect 21968 18470 21980 18522
rect 22032 18470 22044 18522
rect 22096 18470 28734 18522
rect 28786 18470 28798 18522
rect 28850 18470 28862 18522
rect 28914 18470 28926 18522
rect 28978 18470 28990 18522
rect 29042 18470 29048 18522
rect 1104 18448 29048 18470
rect 1578 18068 1584 18080
rect 1539 18040 1584 18068
rect 1578 18028 1584 18040
rect 1636 18028 1642 18080
rect 1104 17978 28888 18000
rect 1104 17926 4423 17978
rect 4475 17926 4487 17978
rect 4539 17926 4551 17978
rect 4603 17926 4615 17978
rect 4667 17926 4679 17978
rect 4731 17926 11369 17978
rect 11421 17926 11433 17978
rect 11485 17926 11497 17978
rect 11549 17926 11561 17978
rect 11613 17926 11625 17978
rect 11677 17926 18315 17978
rect 18367 17926 18379 17978
rect 18431 17926 18443 17978
rect 18495 17926 18507 17978
rect 18559 17926 18571 17978
rect 18623 17926 25261 17978
rect 25313 17926 25325 17978
rect 25377 17926 25389 17978
rect 25441 17926 25453 17978
rect 25505 17926 25517 17978
rect 25569 17926 28888 17978
rect 1104 17904 28888 17926
rect 1578 17660 1584 17672
rect 1539 17632 1584 17660
rect 1578 17620 1584 17632
rect 1636 17620 1642 17672
rect 28350 17660 28356 17672
rect 28311 17632 28356 17660
rect 28350 17620 28356 17632
rect 28408 17620 28414 17672
rect 1104 17434 29048 17456
rect 1104 17382 7896 17434
rect 7948 17382 7960 17434
rect 8012 17382 8024 17434
rect 8076 17382 8088 17434
rect 8140 17382 8152 17434
rect 8204 17382 14842 17434
rect 14894 17382 14906 17434
rect 14958 17382 14970 17434
rect 15022 17382 15034 17434
rect 15086 17382 15098 17434
rect 15150 17382 21788 17434
rect 21840 17382 21852 17434
rect 21904 17382 21916 17434
rect 21968 17382 21980 17434
rect 22032 17382 22044 17434
rect 22096 17382 28734 17434
rect 28786 17382 28798 17434
rect 28850 17382 28862 17434
rect 28914 17382 28926 17434
rect 28978 17382 28990 17434
rect 29042 17382 29048 17434
rect 1104 17360 29048 17382
rect 28350 16980 28356 16992
rect 28311 16952 28356 16980
rect 28350 16940 28356 16952
rect 28408 16940 28414 16992
rect 1104 16890 28888 16912
rect 1104 16838 4423 16890
rect 4475 16838 4487 16890
rect 4539 16838 4551 16890
rect 4603 16838 4615 16890
rect 4667 16838 4679 16890
rect 4731 16838 11369 16890
rect 11421 16838 11433 16890
rect 11485 16838 11497 16890
rect 11549 16838 11561 16890
rect 11613 16838 11625 16890
rect 11677 16838 18315 16890
rect 18367 16838 18379 16890
rect 18431 16838 18443 16890
rect 18495 16838 18507 16890
rect 18559 16838 18571 16890
rect 18623 16838 25261 16890
rect 25313 16838 25325 16890
rect 25377 16838 25389 16890
rect 25441 16838 25453 16890
rect 25505 16838 25517 16890
rect 25569 16838 28888 16890
rect 1104 16816 28888 16838
rect 1104 16346 29048 16368
rect 1104 16294 7896 16346
rect 7948 16294 7960 16346
rect 8012 16294 8024 16346
rect 8076 16294 8088 16346
rect 8140 16294 8152 16346
rect 8204 16294 14842 16346
rect 14894 16294 14906 16346
rect 14958 16294 14970 16346
rect 15022 16294 15034 16346
rect 15086 16294 15098 16346
rect 15150 16294 21788 16346
rect 21840 16294 21852 16346
rect 21904 16294 21916 16346
rect 21968 16294 21980 16346
rect 22032 16294 22044 16346
rect 22096 16294 28734 16346
rect 28786 16294 28798 16346
rect 28850 16294 28862 16346
rect 28914 16294 28926 16346
rect 28978 16294 28990 16346
rect 29042 16294 29048 16346
rect 1104 16272 29048 16294
rect 1578 16028 1584 16040
rect 1539 16000 1584 16028
rect 1578 15988 1584 16000
rect 1636 15988 1642 16040
rect 28350 15892 28356 15904
rect 28311 15864 28356 15892
rect 28350 15852 28356 15864
rect 28408 15852 28414 15904
rect 1104 15802 28888 15824
rect 1104 15750 4423 15802
rect 4475 15750 4487 15802
rect 4539 15750 4551 15802
rect 4603 15750 4615 15802
rect 4667 15750 4679 15802
rect 4731 15750 11369 15802
rect 11421 15750 11433 15802
rect 11485 15750 11497 15802
rect 11549 15750 11561 15802
rect 11613 15750 11625 15802
rect 11677 15750 18315 15802
rect 18367 15750 18379 15802
rect 18431 15750 18443 15802
rect 18495 15750 18507 15802
rect 18559 15750 18571 15802
rect 18623 15750 25261 15802
rect 25313 15750 25325 15802
rect 25377 15750 25389 15802
rect 25441 15750 25453 15802
rect 25505 15750 25517 15802
rect 25569 15750 28888 15802
rect 1104 15728 28888 15750
rect 1578 15484 1584 15496
rect 1539 15456 1584 15484
rect 1578 15444 1584 15456
rect 1636 15444 1642 15496
rect 1104 15258 29048 15280
rect 1104 15206 7896 15258
rect 7948 15206 7960 15258
rect 8012 15206 8024 15258
rect 8076 15206 8088 15258
rect 8140 15206 8152 15258
rect 8204 15206 14842 15258
rect 14894 15206 14906 15258
rect 14958 15206 14970 15258
rect 15022 15206 15034 15258
rect 15086 15206 15098 15258
rect 15150 15206 21788 15258
rect 21840 15206 21852 15258
rect 21904 15206 21916 15258
rect 21968 15206 21980 15258
rect 22032 15206 22044 15258
rect 22096 15206 28734 15258
rect 28786 15206 28798 15258
rect 28850 15206 28862 15258
rect 28914 15206 28926 15258
rect 28978 15206 28990 15258
rect 29042 15206 29048 15258
rect 1104 15184 29048 15206
rect 28350 14872 28356 14884
rect 28311 14844 28356 14872
rect 28350 14832 28356 14844
rect 28408 14832 28414 14884
rect 1104 14714 28888 14736
rect 1104 14662 4423 14714
rect 4475 14662 4487 14714
rect 4539 14662 4551 14714
rect 4603 14662 4615 14714
rect 4667 14662 4679 14714
rect 4731 14662 11369 14714
rect 11421 14662 11433 14714
rect 11485 14662 11497 14714
rect 11549 14662 11561 14714
rect 11613 14662 11625 14714
rect 11677 14662 18315 14714
rect 18367 14662 18379 14714
rect 18431 14662 18443 14714
rect 18495 14662 18507 14714
rect 18559 14662 18571 14714
rect 18623 14662 25261 14714
rect 25313 14662 25325 14714
rect 25377 14662 25389 14714
rect 25441 14662 25453 14714
rect 25505 14662 25517 14714
rect 25569 14662 28888 14714
rect 1104 14640 28888 14662
rect 1578 14396 1584 14408
rect 1539 14368 1584 14396
rect 1578 14356 1584 14368
rect 1636 14356 1642 14408
rect 1104 14170 29048 14192
rect 1104 14118 7896 14170
rect 7948 14118 7960 14170
rect 8012 14118 8024 14170
rect 8076 14118 8088 14170
rect 8140 14118 8152 14170
rect 8204 14118 14842 14170
rect 14894 14118 14906 14170
rect 14958 14118 14970 14170
rect 15022 14118 15034 14170
rect 15086 14118 15098 14170
rect 15150 14118 21788 14170
rect 21840 14118 21852 14170
rect 21904 14118 21916 14170
rect 21968 14118 21980 14170
rect 22032 14118 22044 14170
rect 22096 14118 28734 14170
rect 28786 14118 28798 14170
rect 28850 14118 28862 14170
rect 28914 14118 28926 14170
rect 28978 14118 28990 14170
rect 29042 14118 29048 14170
rect 1104 14096 29048 14118
rect 28350 13716 28356 13728
rect 28311 13688 28356 13716
rect 28350 13676 28356 13688
rect 28408 13676 28414 13728
rect 1104 13626 28888 13648
rect 1104 13574 4423 13626
rect 4475 13574 4487 13626
rect 4539 13574 4551 13626
rect 4603 13574 4615 13626
rect 4667 13574 4679 13626
rect 4731 13574 11369 13626
rect 11421 13574 11433 13626
rect 11485 13574 11497 13626
rect 11549 13574 11561 13626
rect 11613 13574 11625 13626
rect 11677 13574 18315 13626
rect 18367 13574 18379 13626
rect 18431 13574 18443 13626
rect 18495 13574 18507 13626
rect 18559 13574 18571 13626
rect 18623 13574 25261 13626
rect 25313 13574 25325 13626
rect 25377 13574 25389 13626
rect 25441 13574 25453 13626
rect 25505 13574 25517 13626
rect 25569 13574 28888 13626
rect 1104 13552 28888 13574
rect 1578 13308 1584 13320
rect 1539 13280 1584 13308
rect 1578 13268 1584 13280
rect 1636 13268 1642 13320
rect 28350 13308 28356 13320
rect 28311 13280 28356 13308
rect 28350 13268 28356 13280
rect 28408 13268 28414 13320
rect 1104 13082 29048 13104
rect 1104 13030 7896 13082
rect 7948 13030 7960 13082
rect 8012 13030 8024 13082
rect 8076 13030 8088 13082
rect 8140 13030 8152 13082
rect 8204 13030 14842 13082
rect 14894 13030 14906 13082
rect 14958 13030 14970 13082
rect 15022 13030 15034 13082
rect 15086 13030 15098 13082
rect 15150 13030 21788 13082
rect 21840 13030 21852 13082
rect 21904 13030 21916 13082
rect 21968 13030 21980 13082
rect 22032 13030 22044 13082
rect 22096 13030 28734 13082
rect 28786 13030 28798 13082
rect 28850 13030 28862 13082
rect 28914 13030 28926 13082
rect 28978 13030 28990 13082
rect 29042 13030 29048 13082
rect 1104 13008 29048 13030
rect 1104 12538 28888 12560
rect 1104 12486 4423 12538
rect 4475 12486 4487 12538
rect 4539 12486 4551 12538
rect 4603 12486 4615 12538
rect 4667 12486 4679 12538
rect 4731 12486 11369 12538
rect 11421 12486 11433 12538
rect 11485 12486 11497 12538
rect 11549 12486 11561 12538
rect 11613 12486 11625 12538
rect 11677 12486 18315 12538
rect 18367 12486 18379 12538
rect 18431 12486 18443 12538
rect 18495 12486 18507 12538
rect 18559 12486 18571 12538
rect 18623 12486 25261 12538
rect 25313 12486 25325 12538
rect 25377 12486 25389 12538
rect 25441 12486 25453 12538
rect 25505 12486 25517 12538
rect 25569 12486 28888 12538
rect 1104 12464 28888 12486
rect 1578 12220 1584 12232
rect 1539 12192 1584 12220
rect 1578 12180 1584 12192
rect 1636 12180 1642 12232
rect 1104 11994 29048 12016
rect 1104 11942 7896 11994
rect 7948 11942 7960 11994
rect 8012 11942 8024 11994
rect 8076 11942 8088 11994
rect 8140 11942 8152 11994
rect 8204 11942 14842 11994
rect 14894 11942 14906 11994
rect 14958 11942 14970 11994
rect 15022 11942 15034 11994
rect 15086 11942 15098 11994
rect 15150 11942 21788 11994
rect 21840 11942 21852 11994
rect 21904 11942 21916 11994
rect 21968 11942 21980 11994
rect 22032 11942 22044 11994
rect 22096 11942 28734 11994
rect 28786 11942 28798 11994
rect 28850 11942 28862 11994
rect 28914 11942 28926 11994
rect 28978 11942 28990 11994
rect 29042 11942 29048 11994
rect 1104 11920 29048 11942
rect 1578 11540 1584 11552
rect 1539 11512 1584 11540
rect 1578 11500 1584 11512
rect 1636 11500 1642 11552
rect 28350 11540 28356 11552
rect 28311 11512 28356 11540
rect 28350 11500 28356 11512
rect 28408 11500 28414 11552
rect 1104 11450 28888 11472
rect 1104 11398 4423 11450
rect 4475 11398 4487 11450
rect 4539 11398 4551 11450
rect 4603 11398 4615 11450
rect 4667 11398 4679 11450
rect 4731 11398 11369 11450
rect 11421 11398 11433 11450
rect 11485 11398 11497 11450
rect 11549 11398 11561 11450
rect 11613 11398 11625 11450
rect 11677 11398 18315 11450
rect 18367 11398 18379 11450
rect 18431 11398 18443 11450
rect 18495 11398 18507 11450
rect 18559 11398 18571 11450
rect 18623 11398 25261 11450
rect 25313 11398 25325 11450
rect 25377 11398 25389 11450
rect 25441 11398 25453 11450
rect 25505 11398 25517 11450
rect 25569 11398 28888 11450
rect 1104 11376 28888 11398
rect 28350 11132 28356 11144
rect 28311 11104 28356 11132
rect 28350 11092 28356 11104
rect 28408 11092 28414 11144
rect 1104 10906 29048 10928
rect 1104 10854 7896 10906
rect 7948 10854 7960 10906
rect 8012 10854 8024 10906
rect 8076 10854 8088 10906
rect 8140 10854 8152 10906
rect 8204 10854 14842 10906
rect 14894 10854 14906 10906
rect 14958 10854 14970 10906
rect 15022 10854 15034 10906
rect 15086 10854 15098 10906
rect 15150 10854 21788 10906
rect 21840 10854 21852 10906
rect 21904 10854 21916 10906
rect 21968 10854 21980 10906
rect 22032 10854 22044 10906
rect 22096 10854 28734 10906
rect 28786 10854 28798 10906
rect 28850 10854 28862 10906
rect 28914 10854 28926 10906
rect 28978 10854 28990 10906
rect 29042 10854 29048 10906
rect 1104 10832 29048 10854
rect 1104 10362 28888 10384
rect 1104 10310 4423 10362
rect 4475 10310 4487 10362
rect 4539 10310 4551 10362
rect 4603 10310 4615 10362
rect 4667 10310 4679 10362
rect 4731 10310 11369 10362
rect 11421 10310 11433 10362
rect 11485 10310 11497 10362
rect 11549 10310 11561 10362
rect 11613 10310 11625 10362
rect 11677 10310 18315 10362
rect 18367 10310 18379 10362
rect 18431 10310 18443 10362
rect 18495 10310 18507 10362
rect 18559 10310 18571 10362
rect 18623 10310 25261 10362
rect 25313 10310 25325 10362
rect 25377 10310 25389 10362
rect 25441 10310 25453 10362
rect 25505 10310 25517 10362
rect 25569 10310 28888 10362
rect 1104 10288 28888 10310
rect 1578 10044 1584 10056
rect 1539 10016 1584 10044
rect 1578 10004 1584 10016
rect 1636 10004 1642 10056
rect 1104 9818 29048 9840
rect 1104 9766 7896 9818
rect 7948 9766 7960 9818
rect 8012 9766 8024 9818
rect 8076 9766 8088 9818
rect 8140 9766 8152 9818
rect 8204 9766 14842 9818
rect 14894 9766 14906 9818
rect 14958 9766 14970 9818
rect 15022 9766 15034 9818
rect 15086 9766 15098 9818
rect 15150 9766 21788 9818
rect 21840 9766 21852 9818
rect 21904 9766 21916 9818
rect 21968 9766 21980 9818
rect 22032 9766 22044 9818
rect 22096 9766 28734 9818
rect 28786 9766 28798 9818
rect 28850 9766 28862 9818
rect 28914 9766 28926 9818
rect 28978 9766 28990 9818
rect 29042 9766 29048 9818
rect 1104 9744 29048 9766
rect 28350 9432 28356 9444
rect 28311 9404 28356 9432
rect 28350 9392 28356 9404
rect 28408 9392 28414 9444
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 1104 9274 28888 9296
rect 1104 9222 4423 9274
rect 4475 9222 4487 9274
rect 4539 9222 4551 9274
rect 4603 9222 4615 9274
rect 4667 9222 4679 9274
rect 4731 9222 11369 9274
rect 11421 9222 11433 9274
rect 11485 9222 11497 9274
rect 11549 9222 11561 9274
rect 11613 9222 11625 9274
rect 11677 9222 18315 9274
rect 18367 9222 18379 9274
rect 18431 9222 18443 9274
rect 18495 9222 18507 9274
rect 18559 9222 18571 9274
rect 18623 9222 25261 9274
rect 25313 9222 25325 9274
rect 25377 9222 25389 9274
rect 25441 9222 25453 9274
rect 25505 9222 25517 9274
rect 25569 9222 28888 9274
rect 1104 9200 28888 9222
rect 28350 9092 28356 9104
rect 28311 9064 28356 9092
rect 28350 9052 28356 9064
rect 28408 9052 28414 9104
rect 1104 8730 29048 8752
rect 1104 8678 7896 8730
rect 7948 8678 7960 8730
rect 8012 8678 8024 8730
rect 8076 8678 8088 8730
rect 8140 8678 8152 8730
rect 8204 8678 14842 8730
rect 14894 8678 14906 8730
rect 14958 8678 14970 8730
rect 15022 8678 15034 8730
rect 15086 8678 15098 8730
rect 15150 8678 21788 8730
rect 21840 8678 21852 8730
rect 21904 8678 21916 8730
rect 21968 8678 21980 8730
rect 22032 8678 22044 8730
rect 22096 8678 28734 8730
rect 28786 8678 28798 8730
rect 28850 8678 28862 8730
rect 28914 8678 28926 8730
rect 28978 8678 28990 8730
rect 29042 8678 29048 8730
rect 1104 8656 29048 8678
rect 1104 8186 28888 8208
rect 1104 8134 4423 8186
rect 4475 8134 4487 8186
rect 4539 8134 4551 8186
rect 4603 8134 4615 8186
rect 4667 8134 4679 8186
rect 4731 8134 11369 8186
rect 11421 8134 11433 8186
rect 11485 8134 11497 8186
rect 11549 8134 11561 8186
rect 11613 8134 11625 8186
rect 11677 8134 18315 8186
rect 18367 8134 18379 8186
rect 18431 8134 18443 8186
rect 18495 8134 18507 8186
rect 18559 8134 18571 8186
rect 18623 8134 25261 8186
rect 25313 8134 25325 8186
rect 25377 8134 25389 8186
rect 25441 8134 25453 8186
rect 25505 8134 25517 8186
rect 25569 8134 28888 8186
rect 1104 8112 28888 8134
rect 1578 7868 1584 7880
rect 1539 7840 1584 7868
rect 1578 7828 1584 7840
rect 1636 7828 1642 7880
rect 28350 7868 28356 7880
rect 28311 7840 28356 7868
rect 28350 7828 28356 7840
rect 28408 7828 28414 7880
rect 1104 7642 29048 7664
rect 1104 7590 7896 7642
rect 7948 7590 7960 7642
rect 8012 7590 8024 7642
rect 8076 7590 8088 7642
rect 8140 7590 8152 7642
rect 8204 7590 14842 7642
rect 14894 7590 14906 7642
rect 14958 7590 14970 7642
rect 15022 7590 15034 7642
rect 15086 7590 15098 7642
rect 15150 7590 21788 7642
rect 21840 7590 21852 7642
rect 21904 7590 21916 7642
rect 21968 7590 21980 7642
rect 22032 7590 22044 7642
rect 22096 7590 28734 7642
rect 28786 7590 28798 7642
rect 28850 7590 28862 7642
rect 28914 7590 28926 7642
rect 28978 7590 28990 7642
rect 29042 7590 29048 7642
rect 1104 7568 29048 7590
rect 1578 7188 1584 7200
rect 1539 7160 1584 7188
rect 1578 7148 1584 7160
rect 1636 7148 1642 7200
rect 1104 7098 28888 7120
rect 1104 7046 4423 7098
rect 4475 7046 4487 7098
rect 4539 7046 4551 7098
rect 4603 7046 4615 7098
rect 4667 7046 4679 7098
rect 4731 7046 11369 7098
rect 11421 7046 11433 7098
rect 11485 7046 11497 7098
rect 11549 7046 11561 7098
rect 11613 7046 11625 7098
rect 11677 7046 18315 7098
rect 18367 7046 18379 7098
rect 18431 7046 18443 7098
rect 18495 7046 18507 7098
rect 18559 7046 18571 7098
rect 18623 7046 25261 7098
rect 25313 7046 25325 7098
rect 25377 7046 25389 7098
rect 25441 7046 25453 7098
rect 25505 7046 25517 7098
rect 25569 7046 28888 7098
rect 1104 7024 28888 7046
rect 28350 6780 28356 6792
rect 28311 6752 28356 6780
rect 28350 6740 28356 6752
rect 28408 6740 28414 6792
rect 1104 6554 29048 6576
rect 1104 6502 7896 6554
rect 7948 6502 7960 6554
rect 8012 6502 8024 6554
rect 8076 6502 8088 6554
rect 8140 6502 8152 6554
rect 8204 6502 14842 6554
rect 14894 6502 14906 6554
rect 14958 6502 14970 6554
rect 15022 6502 15034 6554
rect 15086 6502 15098 6554
rect 15150 6502 21788 6554
rect 21840 6502 21852 6554
rect 21904 6502 21916 6554
rect 21968 6502 21980 6554
rect 22032 6502 22044 6554
rect 22096 6502 28734 6554
rect 28786 6502 28798 6554
rect 28850 6502 28862 6554
rect 28914 6502 28926 6554
rect 28978 6502 28990 6554
rect 29042 6502 29048 6554
rect 1104 6480 29048 6502
rect 1578 6100 1584 6112
rect 1539 6072 1584 6100
rect 1578 6060 1584 6072
rect 1636 6060 1642 6112
rect 1104 6010 28888 6032
rect 1104 5958 4423 6010
rect 4475 5958 4487 6010
rect 4539 5958 4551 6010
rect 4603 5958 4615 6010
rect 4667 5958 4679 6010
rect 4731 5958 11369 6010
rect 11421 5958 11433 6010
rect 11485 5958 11497 6010
rect 11549 5958 11561 6010
rect 11613 5958 11625 6010
rect 11677 5958 18315 6010
rect 18367 5958 18379 6010
rect 18431 5958 18443 6010
rect 18495 5958 18507 6010
rect 18559 5958 18571 6010
rect 18623 5958 25261 6010
rect 25313 5958 25325 6010
rect 25377 5958 25389 6010
rect 25441 5958 25453 6010
rect 25505 5958 25517 6010
rect 25569 5958 28888 6010
rect 1104 5936 28888 5958
rect 28350 5692 28356 5704
rect 28311 5664 28356 5692
rect 28350 5652 28356 5664
rect 28408 5652 28414 5704
rect 1104 5466 29048 5488
rect 1104 5414 7896 5466
rect 7948 5414 7960 5466
rect 8012 5414 8024 5466
rect 8076 5414 8088 5466
rect 8140 5414 8152 5466
rect 8204 5414 14842 5466
rect 14894 5414 14906 5466
rect 14958 5414 14970 5466
rect 15022 5414 15034 5466
rect 15086 5414 15098 5466
rect 15150 5414 21788 5466
rect 21840 5414 21852 5466
rect 21904 5414 21916 5466
rect 21968 5414 21980 5466
rect 22032 5414 22044 5466
rect 22096 5414 28734 5466
rect 28786 5414 28798 5466
rect 28850 5414 28862 5466
rect 28914 5414 28926 5466
rect 28978 5414 28990 5466
rect 29042 5414 29048 5466
rect 1104 5392 29048 5414
rect 1578 5148 1584 5160
rect 1539 5120 1584 5148
rect 1578 5108 1584 5120
rect 1636 5108 1642 5160
rect 28350 5012 28356 5024
rect 28311 4984 28356 5012
rect 28350 4972 28356 4984
rect 28408 4972 28414 5024
rect 1104 4922 28888 4944
rect 1104 4870 4423 4922
rect 4475 4870 4487 4922
rect 4539 4870 4551 4922
rect 4603 4870 4615 4922
rect 4667 4870 4679 4922
rect 4731 4870 11369 4922
rect 11421 4870 11433 4922
rect 11485 4870 11497 4922
rect 11549 4870 11561 4922
rect 11613 4870 11625 4922
rect 11677 4870 18315 4922
rect 18367 4870 18379 4922
rect 18431 4870 18443 4922
rect 18495 4870 18507 4922
rect 18559 4870 18571 4922
rect 18623 4870 25261 4922
rect 25313 4870 25325 4922
rect 25377 4870 25389 4922
rect 25441 4870 25453 4922
rect 25505 4870 25517 4922
rect 25569 4870 28888 4922
rect 1104 4848 28888 4870
rect 28350 4468 28356 4480
rect 28311 4440 28356 4468
rect 28350 4428 28356 4440
rect 28408 4428 28414 4480
rect 1104 4378 29048 4400
rect 1104 4326 7896 4378
rect 7948 4326 7960 4378
rect 8012 4326 8024 4378
rect 8076 4326 8088 4378
rect 8140 4326 8152 4378
rect 8204 4326 14842 4378
rect 14894 4326 14906 4378
rect 14958 4326 14970 4378
rect 15022 4326 15034 4378
rect 15086 4326 15098 4378
rect 15150 4326 21788 4378
rect 21840 4326 21852 4378
rect 21904 4326 21916 4378
rect 21968 4326 21980 4378
rect 22032 4326 22044 4378
rect 22096 4326 28734 4378
rect 28786 4326 28798 4378
rect 28850 4326 28862 4378
rect 28914 4326 28926 4378
rect 28978 4326 28990 4378
rect 29042 4326 29048 4378
rect 1104 4304 29048 4326
rect 17126 4020 17132 4072
rect 17184 4060 17190 4072
rect 28077 4063 28135 4069
rect 28077 4060 28089 4063
rect 17184 4032 28089 4060
rect 17184 4020 17190 4032
rect 28077 4029 28089 4032
rect 28123 4029 28135 4063
rect 28350 4060 28356 4072
rect 28311 4032 28356 4060
rect 28077 4023 28135 4029
rect 28350 4020 28356 4032
rect 28408 4020 28414 4072
rect 1578 3924 1584 3936
rect 1539 3896 1584 3924
rect 1578 3884 1584 3896
rect 1636 3884 1642 3936
rect 1104 3834 28888 3856
rect 1104 3782 4423 3834
rect 4475 3782 4487 3834
rect 4539 3782 4551 3834
rect 4603 3782 4615 3834
rect 4667 3782 4679 3834
rect 4731 3782 11369 3834
rect 11421 3782 11433 3834
rect 11485 3782 11497 3834
rect 11549 3782 11561 3834
rect 11613 3782 11625 3834
rect 11677 3782 18315 3834
rect 18367 3782 18379 3834
rect 18431 3782 18443 3834
rect 18495 3782 18507 3834
rect 18559 3782 18571 3834
rect 18623 3782 25261 3834
rect 25313 3782 25325 3834
rect 25377 3782 25389 3834
rect 25441 3782 25453 3834
rect 25505 3782 25517 3834
rect 25569 3782 28888 3834
rect 1104 3760 28888 3782
rect 28350 3652 28356 3664
rect 28311 3624 28356 3652
rect 28350 3612 28356 3624
rect 28408 3612 28414 3664
rect 1578 3516 1584 3528
rect 1539 3488 1584 3516
rect 1578 3476 1584 3488
rect 1636 3476 1642 3528
rect 1104 3290 29048 3312
rect 1104 3238 7896 3290
rect 7948 3238 7960 3290
rect 8012 3238 8024 3290
rect 8076 3238 8088 3290
rect 8140 3238 8152 3290
rect 8204 3238 14842 3290
rect 14894 3238 14906 3290
rect 14958 3238 14970 3290
rect 15022 3238 15034 3290
rect 15086 3238 15098 3290
rect 15150 3238 21788 3290
rect 21840 3238 21852 3290
rect 21904 3238 21916 3290
rect 21968 3238 21980 3290
rect 22032 3238 22044 3290
rect 22096 3238 28734 3290
rect 28786 3238 28798 3290
rect 28850 3238 28862 3290
rect 28914 3238 28926 3290
rect 28978 3238 28990 3290
rect 29042 3238 29048 3290
rect 1104 3216 29048 3238
rect 28350 2836 28356 2848
rect 28311 2808 28356 2836
rect 28350 2796 28356 2808
rect 28408 2796 28414 2848
rect 1104 2746 28888 2768
rect 1104 2694 4423 2746
rect 4475 2694 4487 2746
rect 4539 2694 4551 2746
rect 4603 2694 4615 2746
rect 4667 2694 4679 2746
rect 4731 2694 11369 2746
rect 11421 2694 11433 2746
rect 11485 2694 11497 2746
rect 11549 2694 11561 2746
rect 11613 2694 11625 2746
rect 11677 2694 18315 2746
rect 18367 2694 18379 2746
rect 18431 2694 18443 2746
rect 18495 2694 18507 2746
rect 18559 2694 18571 2746
rect 18623 2694 25261 2746
rect 25313 2694 25325 2746
rect 25377 2694 25389 2746
rect 25441 2694 25453 2746
rect 25505 2694 25517 2746
rect 25569 2694 28888 2746
rect 1104 2672 28888 2694
rect 1104 2202 29048 2224
rect 1104 2150 7896 2202
rect 7948 2150 7960 2202
rect 8012 2150 8024 2202
rect 8076 2150 8088 2202
rect 8140 2150 8152 2202
rect 8204 2150 14842 2202
rect 14894 2150 14906 2202
rect 14958 2150 14970 2202
rect 15022 2150 15034 2202
rect 15086 2150 15098 2202
rect 15150 2150 21788 2202
rect 21840 2150 21852 2202
rect 21904 2150 21916 2202
rect 21968 2150 21980 2202
rect 22032 2150 22044 2202
rect 22096 2150 28734 2202
rect 28786 2150 28798 2202
rect 28850 2150 28862 2202
rect 28914 2150 28926 2202
rect 28978 2150 28990 2202
rect 29042 2150 29048 2202
rect 1104 2128 29048 2150
<< via1 >>
rect 12532 31900 12584 31952
rect 14924 31900 14976 31952
rect 13820 31832 13872 31884
rect 16120 31832 16172 31884
rect 12992 31764 13044 31816
rect 16396 31764 16448 31816
rect 9312 31696 9364 31748
rect 13636 31696 13688 31748
rect 14280 31696 14332 31748
rect 19708 31696 19760 31748
rect 4160 31628 4212 31680
rect 6552 31628 6604 31680
rect 7104 31628 7156 31680
rect 8576 31628 8628 31680
rect 14556 31628 14608 31680
rect 7896 31526 7948 31578
rect 7960 31526 8012 31578
rect 8024 31526 8076 31578
rect 8088 31526 8140 31578
rect 8152 31526 8204 31578
rect 14842 31526 14894 31578
rect 14906 31526 14958 31578
rect 14970 31526 15022 31578
rect 15034 31526 15086 31578
rect 15098 31526 15150 31578
rect 21788 31526 21840 31578
rect 21852 31526 21904 31578
rect 21916 31526 21968 31578
rect 21980 31526 22032 31578
rect 22044 31526 22096 31578
rect 28734 31526 28786 31578
rect 28798 31526 28850 31578
rect 28862 31526 28914 31578
rect 28926 31526 28978 31578
rect 28990 31526 29042 31578
rect 5356 31424 5408 31476
rect 11336 31424 11388 31476
rect 13636 31467 13688 31476
rect 13636 31433 13645 31467
rect 13645 31433 13679 31467
rect 13679 31433 13688 31467
rect 13636 31424 13688 31433
rect 14096 31424 14148 31476
rect 4160 31331 4212 31340
rect 4160 31297 4169 31331
rect 4169 31297 4203 31331
rect 4203 31297 4212 31331
rect 4160 31288 4212 31297
rect 5540 31356 5592 31408
rect 5448 31288 5500 31340
rect 6552 31331 6604 31340
rect 6552 31297 6561 31331
rect 6561 31297 6595 31331
rect 6595 31297 6604 31331
rect 6552 31288 6604 31297
rect 14188 31356 14240 31408
rect 14556 31399 14608 31408
rect 14556 31365 14590 31399
rect 14590 31365 14608 31399
rect 14556 31356 14608 31365
rect 17224 31356 17276 31408
rect 2044 31263 2096 31272
rect 2044 31229 2053 31263
rect 2053 31229 2087 31263
rect 2087 31229 2096 31263
rect 2044 31220 2096 31229
rect 6276 31220 6328 31272
rect 9680 31288 9732 31340
rect 10048 31331 10100 31340
rect 10048 31297 10082 31331
rect 10082 31297 10100 31331
rect 10048 31288 10100 31297
rect 12992 31288 13044 31340
rect 15660 31288 15712 31340
rect 16120 31331 16172 31340
rect 16120 31297 16129 31331
rect 16129 31297 16163 31331
rect 16163 31297 16172 31331
rect 16120 31288 16172 31297
rect 16580 31288 16632 31340
rect 9404 31220 9456 31272
rect 9772 31263 9824 31272
rect 9772 31229 9781 31263
rect 9781 31229 9815 31263
rect 9815 31229 9824 31263
rect 9772 31220 9824 31229
rect 3056 31084 3108 31136
rect 3976 31084 4028 31136
rect 6736 31127 6788 31136
rect 6736 31093 6745 31127
rect 6745 31093 6779 31127
rect 6779 31093 6788 31127
rect 6736 31084 6788 31093
rect 8392 31084 8444 31136
rect 10048 31084 10100 31136
rect 11980 31220 12032 31272
rect 13084 31263 13136 31272
rect 13084 31229 13093 31263
rect 13093 31229 13127 31263
rect 13127 31229 13136 31263
rect 13084 31220 13136 31229
rect 17868 31220 17920 31272
rect 21364 31356 21416 31408
rect 20444 31331 20496 31340
rect 19708 31220 19760 31272
rect 20444 31297 20453 31331
rect 20453 31297 20487 31331
rect 20487 31297 20496 31331
rect 20444 31288 20496 31297
rect 20536 31331 20588 31340
rect 20536 31297 20545 31331
rect 20545 31297 20579 31331
rect 20579 31297 20588 31331
rect 20536 31288 20588 31297
rect 20720 31288 20772 31340
rect 21548 31288 21600 31340
rect 23756 31288 23808 31340
rect 24860 31288 24912 31340
rect 27068 31288 27120 31340
rect 28172 31331 28224 31340
rect 28172 31297 28181 31331
rect 28181 31297 28215 31331
rect 28215 31297 28224 31331
rect 28172 31288 28224 31297
rect 12072 31152 12124 31204
rect 17960 31152 18012 31204
rect 11060 31084 11112 31136
rect 11336 31084 11388 31136
rect 13452 31084 13504 31136
rect 13912 31084 13964 31136
rect 15568 31084 15620 31136
rect 18052 31084 18104 31136
rect 18144 31084 18196 31136
rect 20168 31152 20220 31204
rect 19616 31127 19668 31136
rect 19616 31093 19625 31127
rect 19625 31093 19659 31127
rect 19659 31093 19668 31127
rect 19616 31084 19668 31093
rect 19892 31084 19944 31136
rect 4423 30982 4475 31034
rect 4487 30982 4539 31034
rect 4551 30982 4603 31034
rect 4615 30982 4667 31034
rect 4679 30982 4731 31034
rect 11369 30982 11421 31034
rect 11433 30982 11485 31034
rect 11497 30982 11549 31034
rect 11561 30982 11613 31034
rect 11625 30982 11677 31034
rect 18315 30982 18367 31034
rect 18379 30982 18431 31034
rect 18443 30982 18495 31034
rect 18507 30982 18559 31034
rect 18571 30982 18623 31034
rect 25261 30982 25313 31034
rect 25325 30982 25377 31034
rect 25389 30982 25441 31034
rect 25453 30982 25505 31034
rect 25517 30982 25569 31034
rect 7196 30880 7248 30932
rect 8576 30923 8628 30932
rect 8576 30889 8585 30923
rect 8585 30889 8619 30923
rect 8619 30889 8628 30923
rect 8576 30880 8628 30889
rect 9772 30880 9824 30932
rect 4712 30744 4764 30796
rect 5080 30744 5132 30796
rect 11336 30812 11388 30864
rect 12164 30744 12216 30796
rect 12992 30880 13044 30932
rect 14188 30880 14240 30932
rect 20444 30880 20496 30932
rect 21364 30923 21416 30932
rect 21364 30889 21373 30923
rect 21373 30889 21407 30923
rect 21407 30889 21416 30923
rect 21364 30880 21416 30889
rect 27712 30923 27764 30932
rect 27712 30889 27721 30923
rect 27721 30889 27755 30923
rect 27755 30889 27764 30923
rect 27712 30880 27764 30889
rect 28356 30923 28408 30932
rect 28356 30889 28365 30923
rect 28365 30889 28399 30923
rect 28399 30889 28408 30923
rect 28356 30880 28408 30889
rect 13360 30812 13412 30864
rect 14556 30812 14608 30864
rect 16120 30812 16172 30864
rect 18788 30812 18840 30864
rect 13268 30744 13320 30796
rect 14004 30744 14056 30796
rect 15660 30787 15712 30796
rect 15660 30753 15669 30787
rect 15669 30753 15703 30787
rect 15703 30753 15712 30787
rect 15660 30744 15712 30753
rect 16856 30744 16908 30796
rect 19248 30744 19300 30796
rect 19800 30812 19852 30864
rect 2044 30719 2096 30728
rect 2044 30685 2053 30719
rect 2053 30685 2087 30719
rect 2087 30685 2096 30719
rect 2044 30676 2096 30685
rect 2688 30676 2740 30728
rect 6184 30676 6236 30728
rect 6644 30676 6696 30728
rect 9220 30676 9272 30728
rect 9312 30719 9364 30728
rect 9312 30685 9321 30719
rect 9321 30685 9355 30719
rect 9355 30685 9364 30719
rect 9312 30676 9364 30685
rect 10968 30676 11020 30728
rect 4068 30608 4120 30660
rect 4252 30608 4304 30660
rect 4344 30540 4396 30592
rect 4712 30583 4764 30592
rect 4712 30549 4721 30583
rect 4721 30549 4755 30583
rect 4755 30549 4764 30583
rect 4712 30540 4764 30549
rect 7288 30540 7340 30592
rect 7564 30608 7616 30660
rect 7656 30608 7708 30660
rect 10600 30608 10652 30660
rect 15108 30676 15160 30728
rect 15384 30719 15436 30728
rect 15384 30685 15402 30719
rect 15402 30685 15436 30719
rect 15384 30676 15436 30685
rect 13268 30608 13320 30660
rect 10876 30540 10928 30592
rect 13636 30583 13688 30592
rect 13636 30549 13645 30583
rect 13645 30549 13679 30583
rect 13679 30549 13688 30583
rect 13636 30540 13688 30549
rect 14556 30608 14608 30660
rect 17316 30719 17368 30728
rect 17316 30685 17325 30719
rect 17325 30685 17359 30719
rect 17359 30685 17368 30719
rect 17316 30676 17368 30685
rect 17500 30719 17552 30728
rect 17500 30685 17509 30719
rect 17509 30685 17543 30719
rect 17543 30685 17552 30719
rect 17500 30676 17552 30685
rect 16212 30608 16264 30660
rect 14372 30540 14424 30592
rect 16304 30583 16356 30592
rect 16304 30549 16313 30583
rect 16313 30549 16347 30583
rect 16347 30549 16356 30583
rect 16304 30540 16356 30549
rect 16764 30608 16816 30660
rect 19064 30676 19116 30728
rect 19524 30719 19576 30728
rect 19524 30685 19533 30719
rect 19533 30685 19567 30719
rect 19567 30685 19576 30719
rect 20168 30719 20220 30728
rect 19524 30676 19576 30685
rect 20168 30685 20177 30719
rect 20177 30685 20211 30719
rect 20211 30685 20220 30719
rect 20168 30676 20220 30685
rect 20352 30719 20404 30728
rect 20352 30685 20361 30719
rect 20361 30685 20395 30719
rect 20395 30685 20404 30719
rect 20352 30676 20404 30685
rect 19708 30608 19760 30660
rect 16488 30583 16540 30592
rect 16488 30549 16497 30583
rect 16497 30549 16531 30583
rect 16531 30549 16540 30583
rect 16488 30540 16540 30549
rect 17040 30540 17092 30592
rect 20536 30608 20588 30660
rect 20260 30583 20312 30592
rect 20260 30549 20269 30583
rect 20269 30549 20303 30583
rect 20303 30549 20312 30583
rect 20260 30540 20312 30549
rect 7896 30438 7948 30490
rect 7960 30438 8012 30490
rect 8024 30438 8076 30490
rect 8088 30438 8140 30490
rect 8152 30438 8204 30490
rect 14842 30438 14894 30490
rect 14906 30438 14958 30490
rect 14970 30438 15022 30490
rect 15034 30438 15086 30490
rect 15098 30438 15150 30490
rect 21788 30438 21840 30490
rect 21852 30438 21904 30490
rect 21916 30438 21968 30490
rect 21980 30438 22032 30490
rect 22044 30438 22096 30490
rect 28734 30438 28786 30490
rect 28798 30438 28850 30490
rect 28862 30438 28914 30490
rect 28926 30438 28978 30490
rect 28990 30438 29042 30490
rect 2044 30243 2096 30252
rect 2044 30209 2053 30243
rect 2053 30209 2087 30243
rect 2087 30209 2096 30243
rect 2044 30200 2096 30209
rect 3056 30311 3108 30320
rect 3056 30277 3090 30311
rect 3090 30277 3108 30311
rect 3056 30268 3108 30277
rect 4160 30268 4212 30320
rect 3332 30200 3384 30252
rect 5540 30336 5592 30388
rect 8392 30336 8444 30388
rect 10324 30336 10376 30388
rect 10416 30336 10468 30388
rect 11152 30336 11204 30388
rect 12808 30336 12860 30388
rect 14372 30336 14424 30388
rect 2688 30132 2740 30184
rect 3056 29996 3108 30048
rect 6092 30268 6144 30320
rect 6644 30311 6696 30320
rect 6644 30277 6653 30311
rect 6653 30277 6687 30311
rect 6687 30277 6696 30311
rect 6644 30268 6696 30277
rect 7012 30268 7064 30320
rect 12900 30268 12952 30320
rect 14188 30268 14240 30320
rect 14832 30268 14884 30320
rect 5908 30200 5960 30252
rect 6368 30200 6420 30252
rect 6644 30132 6696 30184
rect 7288 30200 7340 30252
rect 9036 30200 9088 30252
rect 10876 30200 10928 30252
rect 12992 30200 13044 30252
rect 14924 30243 14976 30252
rect 14924 30209 14933 30243
rect 14933 30209 14967 30243
rect 14967 30209 14976 30243
rect 14924 30200 14976 30209
rect 15476 30200 15528 30252
rect 15660 30311 15712 30320
rect 15660 30277 15669 30311
rect 15669 30277 15703 30311
rect 15703 30277 15712 30311
rect 16212 30336 16264 30388
rect 16488 30336 16540 30388
rect 17316 30336 17368 30388
rect 17500 30336 17552 30388
rect 17684 30336 17736 30388
rect 15660 30268 15712 30277
rect 19616 30268 19668 30320
rect 7656 30175 7708 30184
rect 7656 30141 7665 30175
rect 7665 30141 7699 30175
rect 7699 30141 7708 30175
rect 7656 30132 7708 30141
rect 9496 30175 9548 30184
rect 9496 30141 9505 30175
rect 9505 30141 9539 30175
rect 9539 30141 9548 30175
rect 9496 30132 9548 30141
rect 11060 30132 11112 30184
rect 11704 30175 11756 30184
rect 11704 30141 11713 30175
rect 11713 30141 11747 30175
rect 11747 30141 11756 30175
rect 11704 30132 11756 30141
rect 6368 29996 6420 30048
rect 6828 30039 6880 30048
rect 6828 30005 6837 30039
rect 6837 30005 6871 30039
rect 6871 30005 6880 30039
rect 6828 29996 6880 30005
rect 8944 29996 8996 30048
rect 10692 29996 10744 30048
rect 10968 29996 11020 30048
rect 13084 30039 13136 30048
rect 13084 30005 13093 30039
rect 13093 30005 13127 30039
rect 13127 30005 13136 30039
rect 13084 29996 13136 30005
rect 17868 30200 17920 30252
rect 18052 30200 18104 30252
rect 19524 30243 19576 30252
rect 17592 30132 17644 30184
rect 15108 30064 15160 30116
rect 15660 30064 15712 30116
rect 17224 30064 17276 30116
rect 15200 29996 15252 30048
rect 16948 30039 17000 30048
rect 16948 30005 16957 30039
rect 16957 30005 16991 30039
rect 16991 30005 17000 30039
rect 16948 29996 17000 30005
rect 17132 29996 17184 30048
rect 17500 29996 17552 30048
rect 18052 29996 18104 30048
rect 18236 30064 18288 30116
rect 18972 29996 19024 30048
rect 19524 30209 19533 30243
rect 19533 30209 19567 30243
rect 19567 30209 19576 30243
rect 19524 30200 19576 30209
rect 28356 30039 28408 30048
rect 28356 30005 28365 30039
rect 28365 30005 28399 30039
rect 28399 30005 28408 30039
rect 28356 29996 28408 30005
rect 4423 29894 4475 29946
rect 4487 29894 4539 29946
rect 4551 29894 4603 29946
rect 4615 29894 4667 29946
rect 4679 29894 4731 29946
rect 11369 29894 11421 29946
rect 11433 29894 11485 29946
rect 11497 29894 11549 29946
rect 11561 29894 11613 29946
rect 11625 29894 11677 29946
rect 18315 29894 18367 29946
rect 18379 29894 18431 29946
rect 18443 29894 18495 29946
rect 18507 29894 18559 29946
rect 18571 29894 18623 29946
rect 25261 29894 25313 29946
rect 25325 29894 25377 29946
rect 25389 29894 25441 29946
rect 25453 29894 25505 29946
rect 25517 29894 25569 29946
rect 3976 29724 4028 29776
rect 4804 29724 4856 29776
rect 6092 29792 6144 29844
rect 6828 29792 6880 29844
rect 9680 29792 9732 29844
rect 13820 29792 13872 29844
rect 6736 29724 6788 29776
rect 7012 29724 7064 29776
rect 7196 29767 7248 29776
rect 7196 29733 7205 29767
rect 7205 29733 7239 29767
rect 7239 29733 7248 29767
rect 7196 29724 7248 29733
rect 10508 29724 10560 29776
rect 2688 29588 2740 29640
rect 2596 29520 2648 29572
rect 5724 29656 5776 29708
rect 6828 29656 6880 29708
rect 7288 29656 7340 29708
rect 10692 29656 10744 29708
rect 5172 29588 5224 29640
rect 8484 29588 8536 29640
rect 9496 29588 9548 29640
rect 1952 29452 2004 29504
rect 3700 29452 3752 29504
rect 4068 29452 4120 29504
rect 6276 29520 6328 29572
rect 7380 29520 7432 29572
rect 10232 29588 10284 29640
rect 9772 29520 9824 29572
rect 7748 29452 7800 29504
rect 8576 29452 8628 29504
rect 10968 29588 11020 29640
rect 10784 29495 10836 29504
rect 10784 29461 10793 29495
rect 10793 29461 10827 29495
rect 10827 29461 10836 29495
rect 10784 29452 10836 29461
rect 11796 29724 11848 29776
rect 13268 29724 13320 29776
rect 13084 29699 13136 29708
rect 13084 29665 13093 29699
rect 13093 29665 13127 29699
rect 13127 29665 13136 29699
rect 13084 29656 13136 29665
rect 11980 29588 12032 29640
rect 14464 29724 14516 29776
rect 14740 29792 14792 29844
rect 15292 29835 15344 29844
rect 15292 29801 15301 29835
rect 15301 29801 15335 29835
rect 15335 29801 15344 29835
rect 15292 29792 15344 29801
rect 15384 29792 15436 29844
rect 15752 29792 15804 29844
rect 17224 29792 17276 29844
rect 15844 29724 15896 29776
rect 15936 29724 15988 29776
rect 17868 29724 17920 29776
rect 18144 29724 18196 29776
rect 18696 29767 18748 29776
rect 18696 29733 18705 29767
rect 18705 29733 18739 29767
rect 18739 29733 18748 29767
rect 18696 29724 18748 29733
rect 14924 29656 14976 29708
rect 15108 29656 15160 29708
rect 15200 29656 15252 29708
rect 15292 29656 15344 29708
rect 15384 29656 15436 29708
rect 20260 29792 20312 29844
rect 14556 29631 14608 29640
rect 14556 29597 14565 29631
rect 14565 29597 14599 29631
rect 14599 29597 14608 29631
rect 14556 29588 14608 29597
rect 14740 29588 14792 29640
rect 16212 29631 16264 29640
rect 12716 29520 12768 29572
rect 13912 29520 13964 29572
rect 15292 29520 15344 29572
rect 16212 29597 16221 29631
rect 16221 29597 16255 29631
rect 16255 29597 16264 29631
rect 16212 29588 16264 29597
rect 16580 29631 16632 29640
rect 16580 29597 16589 29631
rect 16589 29597 16623 29631
rect 16623 29597 16632 29631
rect 16580 29588 16632 29597
rect 16672 29631 16724 29640
rect 16672 29597 16681 29631
rect 16681 29597 16715 29631
rect 16715 29597 16724 29631
rect 16672 29588 16724 29597
rect 17224 29588 17276 29640
rect 18696 29631 18748 29640
rect 18696 29597 18705 29631
rect 18705 29597 18739 29631
rect 18739 29597 18748 29631
rect 18696 29588 18748 29597
rect 18880 29631 18932 29640
rect 18880 29597 18889 29631
rect 18889 29597 18923 29631
rect 18923 29597 18932 29631
rect 18880 29588 18932 29597
rect 28356 29631 28408 29640
rect 28356 29597 28365 29631
rect 28365 29597 28399 29631
rect 28399 29597 28408 29631
rect 28356 29588 28408 29597
rect 16028 29520 16080 29572
rect 17592 29520 17644 29572
rect 17776 29520 17828 29572
rect 19524 29520 19576 29572
rect 20352 29520 20404 29572
rect 13544 29452 13596 29504
rect 14648 29495 14700 29504
rect 14648 29461 14657 29495
rect 14657 29461 14691 29495
rect 14691 29461 14700 29495
rect 17132 29495 17184 29504
rect 14648 29452 14700 29461
rect 17132 29461 17141 29495
rect 17141 29461 17175 29495
rect 17175 29461 17184 29495
rect 17132 29452 17184 29461
rect 17316 29495 17368 29504
rect 17316 29461 17343 29495
rect 17343 29461 17368 29495
rect 17316 29452 17368 29461
rect 18052 29495 18104 29504
rect 18052 29461 18061 29495
rect 18061 29461 18095 29495
rect 18095 29461 18104 29495
rect 18052 29452 18104 29461
rect 7896 29350 7948 29402
rect 7960 29350 8012 29402
rect 8024 29350 8076 29402
rect 8088 29350 8140 29402
rect 8152 29350 8204 29402
rect 14842 29350 14894 29402
rect 14906 29350 14958 29402
rect 14970 29350 15022 29402
rect 15034 29350 15086 29402
rect 15098 29350 15150 29402
rect 21788 29350 21840 29402
rect 21852 29350 21904 29402
rect 21916 29350 21968 29402
rect 21980 29350 22032 29402
rect 22044 29350 22096 29402
rect 28734 29350 28786 29402
rect 28798 29350 28850 29402
rect 28862 29350 28914 29402
rect 28926 29350 28978 29402
rect 28990 29350 29042 29402
rect 2320 29291 2372 29300
rect 2320 29257 2329 29291
rect 2329 29257 2363 29291
rect 2363 29257 2372 29291
rect 2320 29248 2372 29257
rect 3424 29248 3476 29300
rect 6000 29291 6052 29300
rect 2688 29180 2740 29232
rect 1952 29155 2004 29164
rect 1952 29121 1961 29155
rect 1961 29121 1995 29155
rect 1995 29121 2004 29155
rect 1952 29112 2004 29121
rect 2136 29155 2188 29164
rect 2136 29121 2145 29155
rect 2145 29121 2179 29155
rect 2179 29121 2188 29155
rect 2136 29112 2188 29121
rect 3056 29155 3108 29164
rect 3056 29121 3090 29155
rect 3090 29121 3108 29155
rect 5448 29180 5500 29232
rect 6000 29257 6009 29291
rect 6009 29257 6043 29291
rect 6043 29257 6052 29291
rect 6000 29248 6052 29257
rect 6460 29248 6512 29300
rect 7288 29248 7340 29300
rect 7656 29248 7708 29300
rect 11704 29248 11756 29300
rect 12164 29248 12216 29300
rect 12256 29248 12308 29300
rect 12532 29248 12584 29300
rect 12900 29248 12952 29300
rect 14464 29248 14516 29300
rect 9772 29180 9824 29232
rect 11060 29180 11112 29232
rect 12072 29180 12124 29232
rect 12624 29180 12676 29232
rect 14832 29248 14884 29300
rect 15384 29248 15436 29300
rect 16672 29248 16724 29300
rect 3056 29112 3108 29121
rect 5264 29112 5316 29164
rect 5356 29112 5408 29164
rect 2228 28908 2280 28960
rect 6184 29112 6236 29164
rect 7748 29112 7800 29164
rect 8852 29112 8904 29164
rect 9588 29155 9640 29164
rect 9588 29121 9597 29155
rect 9597 29121 9631 29155
rect 9631 29121 9640 29155
rect 9588 29112 9640 29121
rect 9864 29112 9916 29164
rect 11244 29112 11296 29164
rect 12348 29112 12400 29164
rect 15108 29112 15160 29164
rect 15292 29180 15344 29232
rect 18052 29248 18104 29300
rect 6368 29044 6420 29096
rect 7564 29044 7616 29096
rect 11336 29044 11388 29096
rect 11796 29044 11848 29096
rect 14924 29044 14976 29096
rect 7748 28976 7800 29028
rect 8300 28976 8352 29028
rect 8392 28976 8444 29028
rect 10968 28976 11020 29028
rect 12256 28976 12308 29028
rect 3976 28908 4028 28960
rect 10324 28908 10376 28960
rect 11796 28908 11848 28960
rect 11888 28908 11940 28960
rect 15016 28976 15068 29028
rect 12716 28908 12768 28960
rect 15752 28976 15804 29028
rect 16672 29112 16724 29164
rect 16028 29044 16080 29096
rect 16212 29044 16264 29096
rect 17224 29112 17276 29164
rect 17500 29112 17552 29164
rect 17776 29155 17828 29164
rect 17776 29121 17785 29155
rect 17785 29121 17819 29155
rect 17819 29121 17828 29155
rect 17776 29112 17828 29121
rect 16856 29019 16908 29028
rect 15384 28908 15436 28960
rect 16304 28908 16356 28960
rect 16856 28985 16865 29019
rect 16865 28985 16899 29019
rect 16899 28985 16908 29019
rect 16856 28976 16908 28985
rect 17592 29019 17644 29028
rect 17592 28985 17601 29019
rect 17601 28985 17635 29019
rect 17635 28985 17644 29019
rect 17592 28976 17644 28985
rect 17040 28908 17092 28960
rect 18788 28976 18840 29028
rect 4423 28806 4475 28858
rect 4487 28806 4539 28858
rect 4551 28806 4603 28858
rect 4615 28806 4667 28858
rect 4679 28806 4731 28858
rect 11369 28806 11421 28858
rect 11433 28806 11485 28858
rect 11497 28806 11549 28858
rect 11561 28806 11613 28858
rect 11625 28806 11677 28858
rect 18315 28806 18367 28858
rect 18379 28806 18431 28858
rect 18443 28806 18495 28858
rect 18507 28806 18559 28858
rect 18571 28806 18623 28858
rect 25261 28806 25313 28858
rect 25325 28806 25377 28858
rect 25389 28806 25441 28858
rect 25453 28806 25505 28858
rect 25517 28806 25569 28858
rect 5540 28747 5592 28756
rect 5540 28713 5549 28747
rect 5549 28713 5583 28747
rect 5583 28713 5592 28747
rect 5540 28704 5592 28713
rect 6460 28704 6512 28756
rect 9588 28704 9640 28756
rect 12348 28704 12400 28756
rect 13452 28704 13504 28756
rect 6828 28636 6880 28688
rect 8576 28636 8628 28688
rect 9496 28636 9548 28688
rect 12164 28636 12216 28688
rect 12256 28636 12308 28688
rect 14096 28704 14148 28756
rect 15476 28704 15528 28756
rect 16120 28704 16172 28756
rect 18696 28704 18748 28756
rect 9864 28568 9916 28620
rect 13176 28568 13228 28620
rect 2688 28500 2740 28552
rect 5816 28500 5868 28552
rect 9588 28500 9640 28552
rect 9772 28500 9824 28552
rect 13636 28611 13688 28620
rect 13636 28577 13645 28611
rect 13645 28577 13679 28611
rect 13679 28577 13688 28611
rect 13636 28568 13688 28577
rect 14280 28568 14332 28620
rect 14740 28568 14792 28620
rect 14924 28611 14976 28620
rect 14924 28577 14933 28611
rect 14933 28577 14967 28611
rect 14967 28577 14976 28611
rect 14924 28568 14976 28577
rect 16304 28636 16356 28688
rect 18144 28636 18196 28688
rect 15936 28568 15988 28620
rect 16580 28611 16632 28620
rect 16580 28577 16589 28611
rect 16589 28577 16623 28611
rect 16623 28577 16632 28611
rect 16580 28568 16632 28577
rect 4436 28432 4488 28484
rect 5448 28432 5500 28484
rect 7104 28432 7156 28484
rect 4068 28364 4120 28416
rect 8576 28432 8628 28484
rect 8668 28432 8720 28484
rect 12256 28432 12308 28484
rect 12624 28475 12676 28484
rect 12624 28441 12633 28475
rect 12633 28441 12667 28475
rect 12667 28441 12676 28475
rect 12624 28432 12676 28441
rect 7564 28364 7616 28416
rect 10692 28364 10744 28416
rect 10968 28364 11020 28416
rect 12072 28364 12124 28416
rect 13176 28364 13228 28416
rect 13820 28432 13872 28484
rect 14004 28500 14056 28552
rect 14096 28432 14148 28484
rect 13728 28364 13780 28416
rect 15844 28432 15896 28484
rect 16948 28500 17000 28552
rect 17316 28500 17368 28552
rect 17776 28500 17828 28552
rect 7896 28262 7948 28314
rect 7960 28262 8012 28314
rect 8024 28262 8076 28314
rect 8088 28262 8140 28314
rect 8152 28262 8204 28314
rect 14842 28262 14894 28314
rect 14906 28262 14958 28314
rect 14970 28262 15022 28314
rect 15034 28262 15086 28314
rect 15098 28262 15150 28314
rect 21788 28262 21840 28314
rect 21852 28262 21904 28314
rect 21916 28262 21968 28314
rect 21980 28262 22032 28314
rect 22044 28262 22096 28314
rect 28734 28262 28786 28314
rect 28798 28262 28850 28314
rect 28862 28262 28914 28314
rect 28926 28262 28978 28314
rect 28990 28262 29042 28314
rect 5632 28160 5684 28212
rect 5816 28160 5868 28212
rect 8300 28160 8352 28212
rect 12900 28160 12952 28212
rect 12992 28160 13044 28212
rect 13176 28160 13228 28212
rect 15936 28160 15988 28212
rect 4436 28024 4488 28076
rect 5540 28092 5592 28144
rect 4896 28067 4948 28076
rect 4896 28033 4930 28067
rect 4930 28033 4948 28067
rect 4896 28024 4948 28033
rect 5724 28024 5776 28076
rect 7104 28024 7156 28076
rect 8484 28092 8536 28144
rect 9956 28092 10008 28144
rect 7656 28024 7708 28076
rect 14740 28024 14792 28076
rect 15016 28067 15068 28076
rect 15016 28033 15025 28067
rect 15025 28033 15059 28067
rect 15059 28033 15068 28067
rect 15016 28024 15068 28033
rect 15844 28067 15896 28076
rect 6460 27956 6512 28008
rect 3608 27888 3660 27940
rect 2320 27820 2372 27872
rect 4160 27820 4212 27872
rect 7196 27956 7248 28008
rect 11704 27999 11756 28008
rect 11704 27965 11713 27999
rect 11713 27965 11747 27999
rect 11747 27965 11756 27999
rect 11704 27956 11756 27965
rect 14372 27999 14424 28008
rect 14372 27965 14381 27999
rect 14381 27965 14415 27999
rect 14415 27965 14424 27999
rect 14372 27956 14424 27965
rect 15844 28033 15853 28067
rect 15853 28033 15887 28067
rect 15887 28033 15896 28067
rect 15844 28024 15896 28033
rect 15936 28067 15988 28076
rect 15936 28033 15945 28067
rect 15945 28033 15979 28067
rect 15979 28033 15988 28067
rect 15936 28024 15988 28033
rect 7564 27888 7616 27940
rect 12716 27888 12768 27940
rect 15476 27956 15528 28008
rect 16488 27956 16540 28008
rect 15108 27888 15160 27940
rect 16580 27888 16632 27940
rect 6092 27820 6144 27872
rect 6368 27820 6420 27872
rect 8576 27820 8628 27872
rect 12992 27820 13044 27872
rect 13268 27820 13320 27872
rect 13452 27820 13504 27872
rect 13912 27863 13964 27872
rect 13912 27829 13921 27863
rect 13921 27829 13955 27863
rect 13955 27829 13964 27863
rect 13912 27820 13964 27829
rect 14280 27863 14332 27872
rect 14280 27829 14289 27863
rect 14289 27829 14323 27863
rect 14323 27829 14332 27863
rect 14280 27820 14332 27829
rect 15384 27820 15436 27872
rect 16028 27820 16080 27872
rect 18880 27820 18932 27872
rect 28356 27863 28408 27872
rect 28356 27829 28365 27863
rect 28365 27829 28399 27863
rect 28399 27829 28408 27863
rect 28356 27820 28408 27829
rect 4423 27718 4475 27770
rect 4487 27718 4539 27770
rect 4551 27718 4603 27770
rect 4615 27718 4667 27770
rect 4679 27718 4731 27770
rect 11369 27718 11421 27770
rect 11433 27718 11485 27770
rect 11497 27718 11549 27770
rect 11561 27718 11613 27770
rect 11625 27718 11677 27770
rect 18315 27718 18367 27770
rect 18379 27718 18431 27770
rect 18443 27718 18495 27770
rect 18507 27718 18559 27770
rect 18571 27718 18623 27770
rect 25261 27718 25313 27770
rect 25325 27718 25377 27770
rect 25389 27718 25441 27770
rect 25453 27718 25505 27770
rect 25517 27718 25569 27770
rect 4896 27616 4948 27668
rect 3424 27591 3476 27600
rect 3424 27557 3433 27591
rect 3433 27557 3467 27591
rect 3467 27557 3476 27591
rect 3424 27548 3476 27557
rect 2596 27480 2648 27532
rect 5172 27548 5224 27600
rect 6092 27616 6144 27668
rect 7472 27616 7524 27668
rect 12256 27616 12308 27668
rect 12348 27616 12400 27668
rect 15108 27616 15160 27668
rect 15292 27659 15344 27668
rect 15292 27625 15301 27659
rect 15301 27625 15335 27659
rect 15335 27625 15344 27659
rect 15292 27616 15344 27625
rect 5356 27591 5408 27600
rect 5356 27557 5365 27591
rect 5365 27557 5399 27591
rect 5399 27557 5408 27591
rect 5356 27548 5408 27557
rect 11612 27548 11664 27600
rect 3332 27455 3384 27464
rect 3332 27421 3341 27455
rect 3341 27421 3375 27455
rect 3375 27421 3384 27455
rect 3332 27412 3384 27421
rect 4068 27412 4120 27464
rect 4620 27412 4672 27464
rect 5724 27480 5776 27532
rect 11704 27480 11756 27532
rect 11888 27548 11940 27600
rect 14372 27548 14424 27600
rect 14464 27548 14516 27600
rect 14648 27548 14700 27600
rect 15936 27591 15988 27600
rect 15936 27557 15945 27591
rect 15945 27557 15979 27591
rect 15979 27557 15988 27591
rect 15936 27548 15988 27557
rect 16396 27548 16448 27600
rect 5540 27412 5592 27464
rect 6000 27412 6052 27464
rect 8484 27412 8536 27464
rect 9312 27412 9364 27464
rect 10140 27412 10192 27464
rect 10968 27412 11020 27464
rect 12164 27412 12216 27464
rect 13084 27480 13136 27532
rect 13820 27480 13872 27532
rect 12624 27412 12676 27464
rect 13176 27455 13228 27464
rect 13176 27421 13185 27455
rect 13185 27421 13219 27455
rect 13219 27421 13228 27455
rect 13176 27412 13228 27421
rect 13452 27455 13504 27464
rect 13452 27421 13461 27455
rect 13461 27421 13495 27455
rect 13495 27421 13504 27455
rect 13452 27412 13504 27421
rect 3608 27344 3660 27396
rect 3792 27344 3844 27396
rect 4712 27276 4764 27328
rect 6460 27387 6512 27396
rect 6460 27353 6478 27387
rect 6478 27353 6512 27387
rect 6460 27344 6512 27353
rect 6644 27344 6696 27396
rect 7564 27344 7616 27396
rect 8392 27276 8444 27328
rect 8668 27276 8720 27328
rect 11888 27344 11940 27396
rect 9404 27276 9456 27328
rect 12900 27344 12952 27396
rect 14004 27344 14056 27396
rect 15108 27480 15160 27532
rect 15476 27480 15528 27532
rect 15752 27412 15804 27464
rect 16672 27455 16724 27464
rect 12256 27276 12308 27328
rect 12716 27276 12768 27328
rect 12992 27319 13044 27328
rect 12992 27285 13001 27319
rect 13001 27285 13035 27319
rect 13035 27285 13044 27319
rect 12992 27276 13044 27285
rect 13820 27276 13872 27328
rect 15108 27319 15160 27328
rect 15108 27285 15117 27319
rect 15117 27285 15151 27319
rect 15151 27285 15160 27319
rect 15292 27319 15344 27328
rect 15108 27276 15160 27285
rect 15292 27285 15319 27319
rect 15319 27285 15344 27319
rect 15292 27276 15344 27285
rect 15844 27344 15896 27396
rect 15936 27387 15988 27396
rect 15936 27353 15945 27387
rect 15945 27353 15979 27387
rect 15979 27353 15988 27387
rect 16672 27421 16681 27455
rect 16681 27421 16715 27455
rect 16715 27421 16724 27455
rect 16672 27412 16724 27421
rect 16856 27455 16908 27464
rect 16856 27421 16865 27455
rect 16865 27421 16899 27455
rect 16899 27421 16908 27455
rect 16856 27412 16908 27421
rect 28356 27455 28408 27464
rect 28356 27421 28365 27455
rect 28365 27421 28399 27455
rect 28399 27421 28408 27455
rect 28356 27412 28408 27421
rect 15936 27344 15988 27353
rect 7896 27174 7948 27226
rect 7960 27174 8012 27226
rect 8024 27174 8076 27226
rect 8088 27174 8140 27226
rect 8152 27174 8204 27226
rect 14842 27174 14894 27226
rect 14906 27174 14958 27226
rect 14970 27174 15022 27226
rect 15034 27174 15086 27226
rect 15098 27174 15150 27226
rect 21788 27174 21840 27226
rect 21852 27174 21904 27226
rect 21916 27174 21968 27226
rect 21980 27174 22032 27226
rect 22044 27174 22096 27226
rect 28734 27174 28786 27226
rect 28798 27174 28850 27226
rect 28862 27174 28914 27226
rect 28926 27174 28978 27226
rect 28990 27174 29042 27226
rect 2872 27072 2924 27124
rect 3240 27115 3292 27124
rect 3240 27081 3249 27115
rect 3249 27081 3283 27115
rect 3283 27081 3292 27115
rect 3240 27072 3292 27081
rect 6644 27072 6696 27124
rect 8392 27072 8444 27124
rect 5356 27004 5408 27056
rect 7196 27004 7248 27056
rect 9772 27004 9824 27056
rect 10140 27004 10192 27056
rect 12900 27072 12952 27124
rect 13544 27072 13596 27124
rect 1768 26800 1820 26852
rect 2872 26936 2924 26988
rect 3056 26936 3108 26988
rect 3792 26936 3844 26988
rect 3976 26936 4028 26988
rect 4160 26936 4212 26988
rect 6000 26979 6052 26988
rect 6000 26945 6009 26979
rect 6009 26945 6043 26979
rect 6043 26945 6052 26979
rect 6000 26936 6052 26945
rect 6368 26936 6420 26988
rect 8484 26936 8536 26988
rect 8576 26979 8628 26988
rect 8576 26945 8585 26979
rect 8585 26945 8619 26979
rect 8619 26945 8628 26979
rect 8576 26936 8628 26945
rect 8944 26936 8996 26988
rect 6092 26868 6144 26920
rect 8392 26911 8444 26920
rect 3424 26775 3476 26784
rect 3424 26741 3433 26775
rect 3433 26741 3467 26775
rect 3467 26741 3476 26775
rect 3424 26732 3476 26741
rect 4160 26732 4212 26784
rect 6000 26800 6052 26852
rect 6736 26800 6788 26852
rect 8392 26877 8401 26911
rect 8401 26877 8435 26911
rect 8435 26877 8444 26911
rect 8392 26868 8444 26877
rect 9128 26868 9180 26920
rect 10692 26868 10744 26920
rect 10968 26868 11020 26920
rect 13636 27004 13688 27056
rect 14004 27004 14056 27056
rect 14372 27072 14424 27124
rect 15200 27072 15252 27124
rect 15936 27072 15988 27124
rect 17040 27072 17092 27124
rect 11980 26936 12032 26988
rect 13176 26979 13228 26988
rect 9036 26800 9088 26852
rect 8392 26732 8444 26784
rect 10692 26732 10744 26784
rect 12440 26868 12492 26920
rect 12808 26868 12860 26920
rect 13176 26945 13185 26979
rect 13185 26945 13219 26979
rect 13219 26945 13228 26979
rect 13176 26936 13228 26945
rect 14464 26936 14516 26988
rect 14832 26936 14884 26988
rect 14280 26843 14332 26852
rect 14280 26809 14289 26843
rect 14289 26809 14323 26843
rect 14323 26809 14332 26843
rect 14280 26800 14332 26809
rect 14740 26800 14792 26852
rect 15292 26868 15344 26920
rect 16212 26868 16264 26920
rect 15936 26800 15988 26852
rect 12532 26732 12584 26784
rect 14096 26775 14148 26784
rect 14096 26741 14105 26775
rect 14105 26741 14139 26775
rect 14139 26741 14148 26775
rect 14096 26732 14148 26741
rect 4423 26630 4475 26682
rect 4487 26630 4539 26682
rect 4551 26630 4603 26682
rect 4615 26630 4667 26682
rect 4679 26630 4731 26682
rect 11369 26630 11421 26682
rect 11433 26630 11485 26682
rect 11497 26630 11549 26682
rect 11561 26630 11613 26682
rect 11625 26630 11677 26682
rect 18315 26630 18367 26682
rect 18379 26630 18431 26682
rect 18443 26630 18495 26682
rect 18507 26630 18559 26682
rect 18571 26630 18623 26682
rect 25261 26630 25313 26682
rect 25325 26630 25377 26682
rect 25389 26630 25441 26682
rect 25453 26630 25505 26682
rect 25517 26630 25569 26682
rect 3240 26503 3292 26512
rect 3240 26469 3249 26503
rect 3249 26469 3283 26503
rect 3283 26469 3292 26503
rect 3240 26460 3292 26469
rect 4436 26460 4488 26512
rect 1584 26367 1636 26376
rect 1584 26333 1593 26367
rect 1593 26333 1627 26367
rect 1627 26333 1636 26367
rect 1584 26324 1636 26333
rect 2596 26392 2648 26444
rect 4988 26528 5040 26580
rect 5724 26528 5776 26580
rect 6092 26528 6144 26580
rect 6552 26528 6604 26580
rect 7196 26571 7248 26580
rect 5632 26460 5684 26512
rect 6644 26460 6696 26512
rect 2688 26256 2740 26308
rect 3056 26256 3108 26308
rect 3240 26367 3292 26376
rect 3240 26333 3249 26367
rect 3249 26333 3283 26367
rect 3283 26333 3292 26367
rect 3240 26324 3292 26333
rect 3792 26256 3844 26308
rect 2320 26231 2372 26240
rect 2320 26197 2329 26231
rect 2329 26197 2363 26231
rect 2363 26197 2372 26231
rect 2320 26188 2372 26197
rect 3608 26188 3660 26240
rect 4344 26324 4396 26376
rect 6092 26392 6144 26444
rect 7196 26537 7205 26571
rect 7205 26537 7239 26571
rect 7239 26537 7248 26571
rect 7196 26528 7248 26537
rect 7288 26528 7340 26580
rect 8392 26503 8444 26512
rect 8392 26469 8401 26503
rect 8401 26469 8435 26503
rect 8435 26469 8444 26503
rect 8392 26460 8444 26469
rect 8668 26392 8720 26444
rect 6000 26367 6052 26376
rect 6000 26333 6009 26367
rect 6009 26333 6043 26367
rect 6043 26333 6052 26367
rect 6000 26324 6052 26333
rect 6184 26324 6236 26376
rect 6276 26324 6328 26376
rect 7472 26324 7524 26376
rect 7656 26324 7708 26376
rect 8852 26392 8904 26444
rect 9036 26528 9088 26580
rect 9496 26528 9548 26580
rect 10048 26528 10100 26580
rect 10968 26528 11020 26580
rect 12348 26528 12400 26580
rect 12716 26528 12768 26580
rect 13636 26528 13688 26580
rect 14096 26528 14148 26580
rect 18236 26528 18288 26580
rect 10600 26460 10652 26512
rect 13912 26460 13964 26512
rect 15292 26460 15344 26512
rect 9128 26435 9180 26444
rect 9128 26401 9137 26435
rect 9137 26401 9171 26435
rect 9171 26401 9180 26435
rect 9128 26392 9180 26401
rect 10324 26392 10376 26444
rect 10968 26392 11020 26444
rect 11244 26392 11296 26444
rect 11336 26324 11388 26376
rect 6736 26299 6788 26308
rect 6736 26265 6745 26299
rect 6745 26265 6779 26299
rect 6779 26265 6788 26299
rect 8576 26299 8628 26308
rect 6736 26256 6788 26265
rect 8576 26265 8585 26299
rect 8585 26265 8619 26299
rect 8619 26265 8628 26299
rect 8576 26256 8628 26265
rect 8944 26256 8996 26308
rect 6276 26188 6328 26240
rect 7288 26188 7340 26240
rect 9128 26188 9180 26240
rect 11704 26256 11756 26308
rect 9680 26188 9732 26240
rect 10968 26188 11020 26240
rect 12532 26392 12584 26444
rect 13452 26392 13504 26444
rect 13636 26435 13688 26444
rect 13636 26401 13645 26435
rect 13645 26401 13679 26435
rect 13679 26401 13688 26435
rect 13636 26392 13688 26401
rect 12440 26324 12492 26376
rect 16120 26392 16172 26444
rect 12348 26256 12400 26308
rect 13084 26256 13136 26308
rect 13360 26256 13412 26308
rect 14188 26324 14240 26376
rect 14464 26367 14516 26376
rect 14464 26333 14473 26367
rect 14473 26333 14507 26367
rect 14507 26333 14516 26367
rect 14464 26324 14516 26333
rect 17592 26324 17644 26376
rect 13176 26188 13228 26240
rect 14464 26188 14516 26240
rect 15476 26231 15528 26240
rect 15476 26197 15485 26231
rect 15485 26197 15519 26231
rect 15519 26197 15528 26231
rect 15476 26188 15528 26197
rect 7896 26086 7948 26138
rect 7960 26086 8012 26138
rect 8024 26086 8076 26138
rect 8088 26086 8140 26138
rect 8152 26086 8204 26138
rect 14842 26086 14894 26138
rect 14906 26086 14958 26138
rect 14970 26086 15022 26138
rect 15034 26086 15086 26138
rect 15098 26086 15150 26138
rect 21788 26086 21840 26138
rect 21852 26086 21904 26138
rect 21916 26086 21968 26138
rect 21980 26086 22032 26138
rect 22044 26086 22096 26138
rect 28734 26086 28786 26138
rect 28798 26086 28850 26138
rect 28862 26086 28914 26138
rect 28926 26086 28978 26138
rect 28990 26086 29042 26138
rect 1676 26027 1728 26036
rect 1676 25993 1685 26027
rect 1685 25993 1719 26027
rect 1719 25993 1728 26027
rect 1676 25984 1728 25993
rect 4896 25984 4948 26036
rect 4160 25916 4212 25968
rect 5632 25916 5684 25968
rect 6552 25959 6604 25968
rect 6552 25925 6561 25959
rect 6561 25925 6595 25959
rect 6595 25925 6604 25959
rect 6552 25916 6604 25925
rect 3884 25848 3936 25900
rect 5540 25848 5592 25900
rect 6184 25848 6236 25900
rect 6276 25848 6328 25900
rect 8484 25984 8536 26036
rect 10508 26027 10560 26036
rect 10508 25993 10517 26027
rect 10517 25993 10551 26027
rect 10551 25993 10560 26027
rect 10508 25984 10560 25993
rect 10968 26027 11020 26036
rect 10968 25993 10977 26027
rect 10977 25993 11011 26027
rect 11011 25993 11020 26027
rect 10968 25984 11020 25993
rect 11336 25984 11388 26036
rect 12164 25984 12216 26036
rect 9588 25959 9640 25968
rect 9588 25925 9597 25959
rect 9597 25925 9631 25959
rect 9631 25925 9640 25959
rect 9588 25916 9640 25925
rect 11704 25959 11756 25968
rect 11704 25925 11713 25959
rect 11713 25925 11747 25959
rect 11747 25925 11756 25959
rect 11704 25916 11756 25925
rect 20 25780 72 25832
rect 6920 25780 6972 25832
rect 7012 25780 7064 25832
rect 9864 25848 9916 25900
rect 10048 25891 10100 25900
rect 10048 25857 10057 25891
rect 10057 25857 10091 25891
rect 10091 25857 10100 25891
rect 10048 25848 10100 25857
rect 10324 25891 10376 25900
rect 10324 25857 10333 25891
rect 10333 25857 10367 25891
rect 10367 25857 10376 25891
rect 10324 25848 10376 25857
rect 12624 25916 12676 25968
rect 12992 25959 13044 25968
rect 12992 25925 13001 25959
rect 13001 25925 13035 25959
rect 13035 25925 13044 25959
rect 12992 25916 13044 25925
rect 14740 25959 14792 25968
rect 13176 25848 13228 25900
rect 11152 25780 11204 25832
rect 13084 25780 13136 25832
rect 13544 25848 13596 25900
rect 13912 25848 13964 25900
rect 14740 25925 14749 25959
rect 14749 25925 14783 25959
rect 14783 25925 14792 25959
rect 14740 25916 14792 25925
rect 15384 25848 15436 25900
rect 17132 25891 17184 25900
rect 17132 25857 17141 25891
rect 17141 25857 17175 25891
rect 17175 25857 17184 25891
rect 17132 25848 17184 25857
rect 15476 25780 15528 25832
rect 2136 25712 2188 25764
rect 4988 25712 5040 25764
rect 6092 25712 6144 25764
rect 7196 25712 7248 25764
rect 7840 25712 7892 25764
rect 9312 25712 9364 25764
rect 9864 25712 9916 25764
rect 11060 25712 11112 25764
rect 2320 25687 2372 25696
rect 2320 25653 2329 25687
rect 2329 25653 2363 25687
rect 2363 25653 2372 25687
rect 2320 25644 2372 25653
rect 4068 25644 4120 25696
rect 8116 25644 8168 25696
rect 11980 25712 12032 25764
rect 12072 25687 12124 25696
rect 12072 25653 12081 25687
rect 12081 25653 12115 25687
rect 12115 25653 12124 25687
rect 16856 25712 16908 25764
rect 28356 25755 28408 25764
rect 28356 25721 28365 25755
rect 28365 25721 28399 25755
rect 28399 25721 28408 25755
rect 28356 25712 28408 25721
rect 12624 25687 12676 25696
rect 12072 25644 12124 25653
rect 12624 25653 12633 25687
rect 12633 25653 12667 25687
rect 12667 25653 12676 25687
rect 12624 25644 12676 25653
rect 12716 25644 12768 25696
rect 13268 25644 13320 25696
rect 17408 25644 17460 25696
rect 4423 25542 4475 25594
rect 4487 25542 4539 25594
rect 4551 25542 4603 25594
rect 4615 25542 4667 25594
rect 4679 25542 4731 25594
rect 11369 25542 11421 25594
rect 11433 25542 11485 25594
rect 11497 25542 11549 25594
rect 11561 25542 11613 25594
rect 11625 25542 11677 25594
rect 18315 25542 18367 25594
rect 18379 25542 18431 25594
rect 18443 25542 18495 25594
rect 18507 25542 18559 25594
rect 18571 25542 18623 25594
rect 25261 25542 25313 25594
rect 25325 25542 25377 25594
rect 25389 25542 25441 25594
rect 25453 25542 25505 25594
rect 25517 25542 25569 25594
rect 2964 25440 3016 25492
rect 4988 25440 5040 25492
rect 7472 25440 7524 25492
rect 8944 25440 8996 25492
rect 12072 25440 12124 25492
rect 12532 25440 12584 25492
rect 2780 25372 2832 25424
rect 5448 25372 5500 25424
rect 5908 25372 5960 25424
rect 9036 25372 9088 25424
rect 3424 25304 3476 25356
rect 7104 25304 7156 25356
rect 8116 25347 8168 25356
rect 6184 25279 6236 25288
rect 6184 25245 6193 25279
rect 6193 25245 6227 25279
rect 6227 25245 6236 25279
rect 6184 25236 6236 25245
rect 8116 25313 8125 25347
rect 8125 25313 8159 25347
rect 8159 25313 8168 25347
rect 8116 25304 8168 25313
rect 3056 25168 3108 25220
rect 6460 25168 6512 25220
rect 6736 25168 6788 25220
rect 4252 25143 4304 25152
rect 4252 25109 4261 25143
rect 4261 25109 4295 25143
rect 4295 25109 4304 25143
rect 7472 25168 7524 25220
rect 8392 25279 8444 25288
rect 8392 25245 8401 25279
rect 8401 25245 8435 25279
rect 8435 25245 8444 25279
rect 8392 25236 8444 25245
rect 8852 25304 8904 25356
rect 9772 25304 9824 25356
rect 9680 25236 9732 25288
rect 9864 25279 9916 25288
rect 9864 25245 9873 25279
rect 9873 25245 9907 25279
rect 9907 25245 9916 25279
rect 9864 25236 9916 25245
rect 9956 25279 10008 25288
rect 9956 25245 9965 25279
rect 9965 25245 9999 25279
rect 9999 25245 10008 25279
rect 10968 25372 11020 25424
rect 11980 25372 12032 25424
rect 14280 25372 14332 25424
rect 28356 25415 28408 25424
rect 28356 25381 28365 25415
rect 28365 25381 28399 25415
rect 28399 25381 28408 25415
rect 28356 25372 28408 25381
rect 9956 25236 10008 25245
rect 11060 25236 11112 25288
rect 11152 25236 11204 25288
rect 11796 25236 11848 25288
rect 16580 25304 16632 25356
rect 11980 25168 12032 25220
rect 12348 25168 12400 25220
rect 13084 25236 13136 25288
rect 12716 25168 12768 25220
rect 17684 25168 17736 25220
rect 7564 25143 7616 25152
rect 4252 25100 4304 25109
rect 7564 25109 7573 25143
rect 7573 25109 7607 25143
rect 7607 25109 7616 25143
rect 9128 25143 9180 25152
rect 7564 25100 7616 25109
rect 9128 25109 9137 25143
rect 9137 25109 9171 25143
rect 9171 25109 9180 25143
rect 9128 25100 9180 25109
rect 10600 25143 10652 25152
rect 10600 25109 10609 25143
rect 10609 25109 10643 25143
rect 10643 25109 10652 25143
rect 10600 25100 10652 25109
rect 12072 25143 12124 25152
rect 12072 25109 12081 25143
rect 12081 25109 12115 25143
rect 12115 25109 12124 25143
rect 12072 25100 12124 25109
rect 14004 25100 14056 25152
rect 14280 25143 14332 25152
rect 14280 25109 14289 25143
rect 14289 25109 14323 25143
rect 14323 25109 14332 25143
rect 14280 25100 14332 25109
rect 7896 24998 7948 25050
rect 7960 24998 8012 25050
rect 8024 24998 8076 25050
rect 8088 24998 8140 25050
rect 8152 24998 8204 25050
rect 14842 24998 14894 25050
rect 14906 24998 14958 25050
rect 14970 24998 15022 25050
rect 15034 24998 15086 25050
rect 15098 24998 15150 25050
rect 21788 24998 21840 25050
rect 21852 24998 21904 25050
rect 21916 24998 21968 25050
rect 21980 24998 22032 25050
rect 22044 24998 22096 25050
rect 28734 24998 28786 25050
rect 28798 24998 28850 25050
rect 28862 24998 28914 25050
rect 28926 24998 28978 25050
rect 28990 24998 29042 25050
rect 2228 24896 2280 24948
rect 6184 24896 6236 24948
rect 3240 24760 3292 24812
rect 4252 24760 4304 24812
rect 5080 24760 5132 24812
rect 7104 24828 7156 24880
rect 7564 24828 7616 24880
rect 8208 24871 8260 24880
rect 8208 24837 8217 24871
rect 8217 24837 8251 24871
rect 8251 24837 8260 24871
rect 8208 24828 8260 24837
rect 8300 24828 8352 24880
rect 9588 24871 9640 24880
rect 6920 24803 6972 24812
rect 6920 24769 6929 24803
rect 6929 24769 6963 24803
rect 6963 24769 6972 24803
rect 6920 24760 6972 24769
rect 2688 24735 2740 24744
rect 2688 24701 2697 24735
rect 2697 24701 2731 24735
rect 2731 24701 2740 24735
rect 2688 24692 2740 24701
rect 2872 24692 2924 24744
rect 6460 24692 6512 24744
rect 6828 24692 6880 24744
rect 4804 24624 4856 24676
rect 9588 24837 9597 24871
rect 9597 24837 9631 24871
rect 9631 24837 9640 24871
rect 9588 24828 9640 24837
rect 9772 24896 9824 24948
rect 12348 24896 12400 24948
rect 13820 24828 13872 24880
rect 8208 24692 8260 24744
rect 10416 24760 10468 24812
rect 10692 24760 10744 24812
rect 11888 24803 11940 24812
rect 11888 24769 11897 24803
rect 11897 24769 11931 24803
rect 11931 24769 11940 24803
rect 11888 24760 11940 24769
rect 11980 24803 12032 24812
rect 11980 24769 11989 24803
rect 11989 24769 12023 24803
rect 12023 24769 12032 24803
rect 11980 24760 12032 24769
rect 9588 24692 9640 24744
rect 6276 24556 6328 24608
rect 7748 24624 7800 24676
rect 7564 24556 7616 24608
rect 10968 24624 11020 24676
rect 8484 24556 8536 24608
rect 9496 24556 9548 24608
rect 10784 24599 10836 24608
rect 10784 24565 10793 24599
rect 10793 24565 10827 24599
rect 10827 24565 10836 24599
rect 11152 24692 11204 24744
rect 12900 24760 12952 24812
rect 13360 24803 13412 24812
rect 13360 24769 13369 24803
rect 13369 24769 13403 24803
rect 13403 24769 13412 24803
rect 13360 24760 13412 24769
rect 13912 24760 13964 24812
rect 14740 24760 14792 24812
rect 11704 24667 11756 24676
rect 11704 24633 11713 24667
rect 11713 24633 11747 24667
rect 11747 24633 11756 24667
rect 11704 24624 11756 24633
rect 10784 24556 10836 24565
rect 12256 24556 12308 24608
rect 4423 24454 4475 24506
rect 4487 24454 4539 24506
rect 4551 24454 4603 24506
rect 4615 24454 4667 24506
rect 4679 24454 4731 24506
rect 11369 24454 11421 24506
rect 11433 24454 11485 24506
rect 11497 24454 11549 24506
rect 11561 24454 11613 24506
rect 11625 24454 11677 24506
rect 18315 24454 18367 24506
rect 18379 24454 18431 24506
rect 18443 24454 18495 24506
rect 18507 24454 18559 24506
rect 18571 24454 18623 24506
rect 25261 24454 25313 24506
rect 25325 24454 25377 24506
rect 25389 24454 25441 24506
rect 25453 24454 25505 24506
rect 25517 24454 25569 24506
rect 2872 24352 2924 24404
rect 4896 24352 4948 24404
rect 8392 24395 8444 24404
rect 8392 24361 8401 24395
rect 8401 24361 8435 24395
rect 8435 24361 8444 24395
rect 8392 24352 8444 24361
rect 8668 24352 8720 24404
rect 9772 24352 9824 24404
rect 9956 24395 10008 24404
rect 9956 24361 9965 24395
rect 9965 24361 9999 24395
rect 9999 24361 10008 24395
rect 9956 24352 10008 24361
rect 10876 24352 10928 24404
rect 10968 24352 11020 24404
rect 11796 24352 11848 24404
rect 3976 24284 4028 24336
rect 16672 24284 16724 24336
rect 5448 24216 5500 24268
rect 6920 24216 6972 24268
rect 7104 24216 7156 24268
rect 1584 24191 1636 24200
rect 1584 24157 1593 24191
rect 1593 24157 1627 24191
rect 1627 24157 1636 24191
rect 1584 24148 1636 24157
rect 6368 24148 6420 24200
rect 8484 24148 8536 24200
rect 8668 24148 8720 24200
rect 9220 24148 9272 24200
rect 9588 24216 9640 24268
rect 9864 24191 9916 24200
rect 9864 24157 9873 24191
rect 9873 24157 9907 24191
rect 9907 24157 9916 24191
rect 9864 24148 9916 24157
rect 12072 24216 12124 24268
rect 10784 24191 10836 24200
rect 10784 24157 10793 24191
rect 10793 24157 10827 24191
rect 10827 24157 10836 24191
rect 10784 24148 10836 24157
rect 28356 24191 28408 24200
rect 28356 24157 28365 24191
rect 28365 24157 28399 24191
rect 28399 24157 28408 24191
rect 28356 24148 28408 24157
rect 7564 24080 7616 24132
rect 7656 24080 7708 24132
rect 10416 24080 10468 24132
rect 11152 24080 11204 24132
rect 6460 24055 6512 24064
rect 6460 24021 6469 24055
rect 6469 24021 6503 24055
rect 6503 24021 6512 24055
rect 6460 24012 6512 24021
rect 7472 24012 7524 24064
rect 7896 23910 7948 23962
rect 7960 23910 8012 23962
rect 8024 23910 8076 23962
rect 8088 23910 8140 23962
rect 8152 23910 8204 23962
rect 14842 23910 14894 23962
rect 14906 23910 14958 23962
rect 14970 23910 15022 23962
rect 15034 23910 15086 23962
rect 15098 23910 15150 23962
rect 21788 23910 21840 23962
rect 21852 23910 21904 23962
rect 21916 23910 21968 23962
rect 21980 23910 22032 23962
rect 22044 23910 22096 23962
rect 28734 23910 28786 23962
rect 28798 23910 28850 23962
rect 28862 23910 28914 23962
rect 28926 23910 28978 23962
rect 28990 23910 29042 23962
rect 5448 23808 5500 23860
rect 6920 23851 6972 23860
rect 6920 23817 6929 23851
rect 6929 23817 6963 23851
rect 6963 23817 6972 23851
rect 6920 23808 6972 23817
rect 7380 23808 7432 23860
rect 5080 23740 5132 23792
rect 10416 23740 10468 23792
rect 8576 23672 8628 23724
rect 14280 23808 14332 23860
rect 6920 23604 6972 23656
rect 8668 23647 8720 23656
rect 8668 23613 8677 23647
rect 8677 23613 8711 23647
rect 8711 23613 8720 23647
rect 8668 23604 8720 23613
rect 9588 23604 9640 23656
rect 1584 23511 1636 23520
rect 1584 23477 1593 23511
rect 1593 23477 1627 23511
rect 1627 23477 1636 23511
rect 1584 23468 1636 23477
rect 6460 23468 6512 23520
rect 13912 23468 13964 23520
rect 4423 23366 4475 23418
rect 4487 23366 4539 23418
rect 4551 23366 4603 23418
rect 4615 23366 4667 23418
rect 4679 23366 4731 23418
rect 11369 23366 11421 23418
rect 11433 23366 11485 23418
rect 11497 23366 11549 23418
rect 11561 23366 11613 23418
rect 11625 23366 11677 23418
rect 18315 23366 18367 23418
rect 18379 23366 18431 23418
rect 18443 23366 18495 23418
rect 18507 23366 18559 23418
rect 18571 23366 18623 23418
rect 25261 23366 25313 23418
rect 25325 23366 25377 23418
rect 25389 23366 25441 23418
rect 25453 23366 25505 23418
rect 25517 23366 25569 23418
rect 9220 23264 9272 23316
rect 28356 23103 28408 23112
rect 28356 23069 28365 23103
rect 28365 23069 28399 23103
rect 28399 23069 28408 23103
rect 28356 23060 28408 23069
rect 7896 22822 7948 22874
rect 7960 22822 8012 22874
rect 8024 22822 8076 22874
rect 8088 22822 8140 22874
rect 8152 22822 8204 22874
rect 14842 22822 14894 22874
rect 14906 22822 14958 22874
rect 14970 22822 15022 22874
rect 15034 22822 15086 22874
rect 15098 22822 15150 22874
rect 21788 22822 21840 22874
rect 21852 22822 21904 22874
rect 21916 22822 21968 22874
rect 21980 22822 22032 22874
rect 22044 22822 22096 22874
rect 28734 22822 28786 22874
rect 28798 22822 28850 22874
rect 28862 22822 28914 22874
rect 28926 22822 28978 22874
rect 28990 22822 29042 22874
rect 1584 22423 1636 22432
rect 1584 22389 1593 22423
rect 1593 22389 1627 22423
rect 1627 22389 1636 22423
rect 1584 22380 1636 22389
rect 4423 22278 4475 22330
rect 4487 22278 4539 22330
rect 4551 22278 4603 22330
rect 4615 22278 4667 22330
rect 4679 22278 4731 22330
rect 11369 22278 11421 22330
rect 11433 22278 11485 22330
rect 11497 22278 11549 22330
rect 11561 22278 11613 22330
rect 11625 22278 11677 22330
rect 18315 22278 18367 22330
rect 18379 22278 18431 22330
rect 18443 22278 18495 22330
rect 18507 22278 18559 22330
rect 18571 22278 18623 22330
rect 25261 22278 25313 22330
rect 25325 22278 25377 22330
rect 25389 22278 25441 22330
rect 25453 22278 25505 22330
rect 25517 22278 25569 22330
rect 28356 22015 28408 22024
rect 28356 21981 28365 22015
rect 28365 21981 28399 22015
rect 28399 21981 28408 22015
rect 28356 21972 28408 21981
rect 7896 21734 7948 21786
rect 7960 21734 8012 21786
rect 8024 21734 8076 21786
rect 8088 21734 8140 21786
rect 8152 21734 8204 21786
rect 14842 21734 14894 21786
rect 14906 21734 14958 21786
rect 14970 21734 15022 21786
rect 15034 21734 15086 21786
rect 15098 21734 15150 21786
rect 21788 21734 21840 21786
rect 21852 21734 21904 21786
rect 21916 21734 21968 21786
rect 21980 21734 22032 21786
rect 22044 21734 22096 21786
rect 28734 21734 28786 21786
rect 28798 21734 28850 21786
rect 28862 21734 28914 21786
rect 28926 21734 28978 21786
rect 28990 21734 29042 21786
rect 1584 21471 1636 21480
rect 1584 21437 1593 21471
rect 1593 21437 1627 21471
rect 1627 21437 1636 21471
rect 1584 21428 1636 21437
rect 28356 21335 28408 21344
rect 28356 21301 28365 21335
rect 28365 21301 28399 21335
rect 28399 21301 28408 21335
rect 28356 21292 28408 21301
rect 4423 21190 4475 21242
rect 4487 21190 4539 21242
rect 4551 21190 4603 21242
rect 4615 21190 4667 21242
rect 4679 21190 4731 21242
rect 11369 21190 11421 21242
rect 11433 21190 11485 21242
rect 11497 21190 11549 21242
rect 11561 21190 11613 21242
rect 11625 21190 11677 21242
rect 18315 21190 18367 21242
rect 18379 21190 18431 21242
rect 18443 21190 18495 21242
rect 18507 21190 18559 21242
rect 18571 21190 18623 21242
rect 25261 21190 25313 21242
rect 25325 21190 25377 21242
rect 25389 21190 25441 21242
rect 25453 21190 25505 21242
rect 25517 21190 25569 21242
rect 7896 20646 7948 20698
rect 7960 20646 8012 20698
rect 8024 20646 8076 20698
rect 8088 20646 8140 20698
rect 8152 20646 8204 20698
rect 14842 20646 14894 20698
rect 14906 20646 14958 20698
rect 14970 20646 15022 20698
rect 15034 20646 15086 20698
rect 15098 20646 15150 20698
rect 21788 20646 21840 20698
rect 21852 20646 21904 20698
rect 21916 20646 21968 20698
rect 21980 20646 22032 20698
rect 22044 20646 22096 20698
rect 28734 20646 28786 20698
rect 28798 20646 28850 20698
rect 28862 20646 28914 20698
rect 28926 20646 28978 20698
rect 28990 20646 29042 20698
rect 1584 20247 1636 20256
rect 1584 20213 1593 20247
rect 1593 20213 1627 20247
rect 1627 20213 1636 20247
rect 1584 20204 1636 20213
rect 4423 20102 4475 20154
rect 4487 20102 4539 20154
rect 4551 20102 4603 20154
rect 4615 20102 4667 20154
rect 4679 20102 4731 20154
rect 11369 20102 11421 20154
rect 11433 20102 11485 20154
rect 11497 20102 11549 20154
rect 11561 20102 11613 20154
rect 11625 20102 11677 20154
rect 18315 20102 18367 20154
rect 18379 20102 18431 20154
rect 18443 20102 18495 20154
rect 18507 20102 18559 20154
rect 18571 20102 18623 20154
rect 25261 20102 25313 20154
rect 25325 20102 25377 20154
rect 25389 20102 25441 20154
rect 25453 20102 25505 20154
rect 25517 20102 25569 20154
rect 28356 19975 28408 19984
rect 28356 19941 28365 19975
rect 28365 19941 28399 19975
rect 28399 19941 28408 19975
rect 28356 19932 28408 19941
rect 1584 19839 1636 19848
rect 1584 19805 1593 19839
rect 1593 19805 1627 19839
rect 1627 19805 1636 19839
rect 1584 19796 1636 19805
rect 7896 19558 7948 19610
rect 7960 19558 8012 19610
rect 8024 19558 8076 19610
rect 8088 19558 8140 19610
rect 8152 19558 8204 19610
rect 14842 19558 14894 19610
rect 14906 19558 14958 19610
rect 14970 19558 15022 19610
rect 15034 19558 15086 19610
rect 15098 19558 15150 19610
rect 21788 19558 21840 19610
rect 21852 19558 21904 19610
rect 21916 19558 21968 19610
rect 21980 19558 22032 19610
rect 22044 19558 22096 19610
rect 28734 19558 28786 19610
rect 28798 19558 28850 19610
rect 28862 19558 28914 19610
rect 28926 19558 28978 19610
rect 28990 19558 29042 19610
rect 28356 19159 28408 19168
rect 28356 19125 28365 19159
rect 28365 19125 28399 19159
rect 28399 19125 28408 19159
rect 28356 19116 28408 19125
rect 4423 19014 4475 19066
rect 4487 19014 4539 19066
rect 4551 19014 4603 19066
rect 4615 19014 4667 19066
rect 4679 19014 4731 19066
rect 11369 19014 11421 19066
rect 11433 19014 11485 19066
rect 11497 19014 11549 19066
rect 11561 19014 11613 19066
rect 11625 19014 11677 19066
rect 18315 19014 18367 19066
rect 18379 19014 18431 19066
rect 18443 19014 18495 19066
rect 18507 19014 18559 19066
rect 18571 19014 18623 19066
rect 25261 19014 25313 19066
rect 25325 19014 25377 19066
rect 25389 19014 25441 19066
rect 25453 19014 25505 19066
rect 25517 19014 25569 19066
rect 7896 18470 7948 18522
rect 7960 18470 8012 18522
rect 8024 18470 8076 18522
rect 8088 18470 8140 18522
rect 8152 18470 8204 18522
rect 14842 18470 14894 18522
rect 14906 18470 14958 18522
rect 14970 18470 15022 18522
rect 15034 18470 15086 18522
rect 15098 18470 15150 18522
rect 21788 18470 21840 18522
rect 21852 18470 21904 18522
rect 21916 18470 21968 18522
rect 21980 18470 22032 18522
rect 22044 18470 22096 18522
rect 28734 18470 28786 18522
rect 28798 18470 28850 18522
rect 28862 18470 28914 18522
rect 28926 18470 28978 18522
rect 28990 18470 29042 18522
rect 1584 18071 1636 18080
rect 1584 18037 1593 18071
rect 1593 18037 1627 18071
rect 1627 18037 1636 18071
rect 1584 18028 1636 18037
rect 4423 17926 4475 17978
rect 4487 17926 4539 17978
rect 4551 17926 4603 17978
rect 4615 17926 4667 17978
rect 4679 17926 4731 17978
rect 11369 17926 11421 17978
rect 11433 17926 11485 17978
rect 11497 17926 11549 17978
rect 11561 17926 11613 17978
rect 11625 17926 11677 17978
rect 18315 17926 18367 17978
rect 18379 17926 18431 17978
rect 18443 17926 18495 17978
rect 18507 17926 18559 17978
rect 18571 17926 18623 17978
rect 25261 17926 25313 17978
rect 25325 17926 25377 17978
rect 25389 17926 25441 17978
rect 25453 17926 25505 17978
rect 25517 17926 25569 17978
rect 1584 17663 1636 17672
rect 1584 17629 1593 17663
rect 1593 17629 1627 17663
rect 1627 17629 1636 17663
rect 1584 17620 1636 17629
rect 28356 17663 28408 17672
rect 28356 17629 28365 17663
rect 28365 17629 28399 17663
rect 28399 17629 28408 17663
rect 28356 17620 28408 17629
rect 7896 17382 7948 17434
rect 7960 17382 8012 17434
rect 8024 17382 8076 17434
rect 8088 17382 8140 17434
rect 8152 17382 8204 17434
rect 14842 17382 14894 17434
rect 14906 17382 14958 17434
rect 14970 17382 15022 17434
rect 15034 17382 15086 17434
rect 15098 17382 15150 17434
rect 21788 17382 21840 17434
rect 21852 17382 21904 17434
rect 21916 17382 21968 17434
rect 21980 17382 22032 17434
rect 22044 17382 22096 17434
rect 28734 17382 28786 17434
rect 28798 17382 28850 17434
rect 28862 17382 28914 17434
rect 28926 17382 28978 17434
rect 28990 17382 29042 17434
rect 28356 16983 28408 16992
rect 28356 16949 28365 16983
rect 28365 16949 28399 16983
rect 28399 16949 28408 16983
rect 28356 16940 28408 16949
rect 4423 16838 4475 16890
rect 4487 16838 4539 16890
rect 4551 16838 4603 16890
rect 4615 16838 4667 16890
rect 4679 16838 4731 16890
rect 11369 16838 11421 16890
rect 11433 16838 11485 16890
rect 11497 16838 11549 16890
rect 11561 16838 11613 16890
rect 11625 16838 11677 16890
rect 18315 16838 18367 16890
rect 18379 16838 18431 16890
rect 18443 16838 18495 16890
rect 18507 16838 18559 16890
rect 18571 16838 18623 16890
rect 25261 16838 25313 16890
rect 25325 16838 25377 16890
rect 25389 16838 25441 16890
rect 25453 16838 25505 16890
rect 25517 16838 25569 16890
rect 7896 16294 7948 16346
rect 7960 16294 8012 16346
rect 8024 16294 8076 16346
rect 8088 16294 8140 16346
rect 8152 16294 8204 16346
rect 14842 16294 14894 16346
rect 14906 16294 14958 16346
rect 14970 16294 15022 16346
rect 15034 16294 15086 16346
rect 15098 16294 15150 16346
rect 21788 16294 21840 16346
rect 21852 16294 21904 16346
rect 21916 16294 21968 16346
rect 21980 16294 22032 16346
rect 22044 16294 22096 16346
rect 28734 16294 28786 16346
rect 28798 16294 28850 16346
rect 28862 16294 28914 16346
rect 28926 16294 28978 16346
rect 28990 16294 29042 16346
rect 1584 16031 1636 16040
rect 1584 15997 1593 16031
rect 1593 15997 1627 16031
rect 1627 15997 1636 16031
rect 1584 15988 1636 15997
rect 28356 15895 28408 15904
rect 28356 15861 28365 15895
rect 28365 15861 28399 15895
rect 28399 15861 28408 15895
rect 28356 15852 28408 15861
rect 4423 15750 4475 15802
rect 4487 15750 4539 15802
rect 4551 15750 4603 15802
rect 4615 15750 4667 15802
rect 4679 15750 4731 15802
rect 11369 15750 11421 15802
rect 11433 15750 11485 15802
rect 11497 15750 11549 15802
rect 11561 15750 11613 15802
rect 11625 15750 11677 15802
rect 18315 15750 18367 15802
rect 18379 15750 18431 15802
rect 18443 15750 18495 15802
rect 18507 15750 18559 15802
rect 18571 15750 18623 15802
rect 25261 15750 25313 15802
rect 25325 15750 25377 15802
rect 25389 15750 25441 15802
rect 25453 15750 25505 15802
rect 25517 15750 25569 15802
rect 1584 15487 1636 15496
rect 1584 15453 1593 15487
rect 1593 15453 1627 15487
rect 1627 15453 1636 15487
rect 1584 15444 1636 15453
rect 7896 15206 7948 15258
rect 7960 15206 8012 15258
rect 8024 15206 8076 15258
rect 8088 15206 8140 15258
rect 8152 15206 8204 15258
rect 14842 15206 14894 15258
rect 14906 15206 14958 15258
rect 14970 15206 15022 15258
rect 15034 15206 15086 15258
rect 15098 15206 15150 15258
rect 21788 15206 21840 15258
rect 21852 15206 21904 15258
rect 21916 15206 21968 15258
rect 21980 15206 22032 15258
rect 22044 15206 22096 15258
rect 28734 15206 28786 15258
rect 28798 15206 28850 15258
rect 28862 15206 28914 15258
rect 28926 15206 28978 15258
rect 28990 15206 29042 15258
rect 28356 14875 28408 14884
rect 28356 14841 28365 14875
rect 28365 14841 28399 14875
rect 28399 14841 28408 14875
rect 28356 14832 28408 14841
rect 4423 14662 4475 14714
rect 4487 14662 4539 14714
rect 4551 14662 4603 14714
rect 4615 14662 4667 14714
rect 4679 14662 4731 14714
rect 11369 14662 11421 14714
rect 11433 14662 11485 14714
rect 11497 14662 11549 14714
rect 11561 14662 11613 14714
rect 11625 14662 11677 14714
rect 18315 14662 18367 14714
rect 18379 14662 18431 14714
rect 18443 14662 18495 14714
rect 18507 14662 18559 14714
rect 18571 14662 18623 14714
rect 25261 14662 25313 14714
rect 25325 14662 25377 14714
rect 25389 14662 25441 14714
rect 25453 14662 25505 14714
rect 25517 14662 25569 14714
rect 1584 14399 1636 14408
rect 1584 14365 1593 14399
rect 1593 14365 1627 14399
rect 1627 14365 1636 14399
rect 1584 14356 1636 14365
rect 7896 14118 7948 14170
rect 7960 14118 8012 14170
rect 8024 14118 8076 14170
rect 8088 14118 8140 14170
rect 8152 14118 8204 14170
rect 14842 14118 14894 14170
rect 14906 14118 14958 14170
rect 14970 14118 15022 14170
rect 15034 14118 15086 14170
rect 15098 14118 15150 14170
rect 21788 14118 21840 14170
rect 21852 14118 21904 14170
rect 21916 14118 21968 14170
rect 21980 14118 22032 14170
rect 22044 14118 22096 14170
rect 28734 14118 28786 14170
rect 28798 14118 28850 14170
rect 28862 14118 28914 14170
rect 28926 14118 28978 14170
rect 28990 14118 29042 14170
rect 28356 13719 28408 13728
rect 28356 13685 28365 13719
rect 28365 13685 28399 13719
rect 28399 13685 28408 13719
rect 28356 13676 28408 13685
rect 4423 13574 4475 13626
rect 4487 13574 4539 13626
rect 4551 13574 4603 13626
rect 4615 13574 4667 13626
rect 4679 13574 4731 13626
rect 11369 13574 11421 13626
rect 11433 13574 11485 13626
rect 11497 13574 11549 13626
rect 11561 13574 11613 13626
rect 11625 13574 11677 13626
rect 18315 13574 18367 13626
rect 18379 13574 18431 13626
rect 18443 13574 18495 13626
rect 18507 13574 18559 13626
rect 18571 13574 18623 13626
rect 25261 13574 25313 13626
rect 25325 13574 25377 13626
rect 25389 13574 25441 13626
rect 25453 13574 25505 13626
rect 25517 13574 25569 13626
rect 1584 13311 1636 13320
rect 1584 13277 1593 13311
rect 1593 13277 1627 13311
rect 1627 13277 1636 13311
rect 1584 13268 1636 13277
rect 28356 13311 28408 13320
rect 28356 13277 28365 13311
rect 28365 13277 28399 13311
rect 28399 13277 28408 13311
rect 28356 13268 28408 13277
rect 7896 13030 7948 13082
rect 7960 13030 8012 13082
rect 8024 13030 8076 13082
rect 8088 13030 8140 13082
rect 8152 13030 8204 13082
rect 14842 13030 14894 13082
rect 14906 13030 14958 13082
rect 14970 13030 15022 13082
rect 15034 13030 15086 13082
rect 15098 13030 15150 13082
rect 21788 13030 21840 13082
rect 21852 13030 21904 13082
rect 21916 13030 21968 13082
rect 21980 13030 22032 13082
rect 22044 13030 22096 13082
rect 28734 13030 28786 13082
rect 28798 13030 28850 13082
rect 28862 13030 28914 13082
rect 28926 13030 28978 13082
rect 28990 13030 29042 13082
rect 4423 12486 4475 12538
rect 4487 12486 4539 12538
rect 4551 12486 4603 12538
rect 4615 12486 4667 12538
rect 4679 12486 4731 12538
rect 11369 12486 11421 12538
rect 11433 12486 11485 12538
rect 11497 12486 11549 12538
rect 11561 12486 11613 12538
rect 11625 12486 11677 12538
rect 18315 12486 18367 12538
rect 18379 12486 18431 12538
rect 18443 12486 18495 12538
rect 18507 12486 18559 12538
rect 18571 12486 18623 12538
rect 25261 12486 25313 12538
rect 25325 12486 25377 12538
rect 25389 12486 25441 12538
rect 25453 12486 25505 12538
rect 25517 12486 25569 12538
rect 1584 12223 1636 12232
rect 1584 12189 1593 12223
rect 1593 12189 1627 12223
rect 1627 12189 1636 12223
rect 1584 12180 1636 12189
rect 7896 11942 7948 11994
rect 7960 11942 8012 11994
rect 8024 11942 8076 11994
rect 8088 11942 8140 11994
rect 8152 11942 8204 11994
rect 14842 11942 14894 11994
rect 14906 11942 14958 11994
rect 14970 11942 15022 11994
rect 15034 11942 15086 11994
rect 15098 11942 15150 11994
rect 21788 11942 21840 11994
rect 21852 11942 21904 11994
rect 21916 11942 21968 11994
rect 21980 11942 22032 11994
rect 22044 11942 22096 11994
rect 28734 11942 28786 11994
rect 28798 11942 28850 11994
rect 28862 11942 28914 11994
rect 28926 11942 28978 11994
rect 28990 11942 29042 11994
rect 1584 11543 1636 11552
rect 1584 11509 1593 11543
rect 1593 11509 1627 11543
rect 1627 11509 1636 11543
rect 1584 11500 1636 11509
rect 28356 11543 28408 11552
rect 28356 11509 28365 11543
rect 28365 11509 28399 11543
rect 28399 11509 28408 11543
rect 28356 11500 28408 11509
rect 4423 11398 4475 11450
rect 4487 11398 4539 11450
rect 4551 11398 4603 11450
rect 4615 11398 4667 11450
rect 4679 11398 4731 11450
rect 11369 11398 11421 11450
rect 11433 11398 11485 11450
rect 11497 11398 11549 11450
rect 11561 11398 11613 11450
rect 11625 11398 11677 11450
rect 18315 11398 18367 11450
rect 18379 11398 18431 11450
rect 18443 11398 18495 11450
rect 18507 11398 18559 11450
rect 18571 11398 18623 11450
rect 25261 11398 25313 11450
rect 25325 11398 25377 11450
rect 25389 11398 25441 11450
rect 25453 11398 25505 11450
rect 25517 11398 25569 11450
rect 28356 11135 28408 11144
rect 28356 11101 28365 11135
rect 28365 11101 28399 11135
rect 28399 11101 28408 11135
rect 28356 11092 28408 11101
rect 7896 10854 7948 10906
rect 7960 10854 8012 10906
rect 8024 10854 8076 10906
rect 8088 10854 8140 10906
rect 8152 10854 8204 10906
rect 14842 10854 14894 10906
rect 14906 10854 14958 10906
rect 14970 10854 15022 10906
rect 15034 10854 15086 10906
rect 15098 10854 15150 10906
rect 21788 10854 21840 10906
rect 21852 10854 21904 10906
rect 21916 10854 21968 10906
rect 21980 10854 22032 10906
rect 22044 10854 22096 10906
rect 28734 10854 28786 10906
rect 28798 10854 28850 10906
rect 28862 10854 28914 10906
rect 28926 10854 28978 10906
rect 28990 10854 29042 10906
rect 4423 10310 4475 10362
rect 4487 10310 4539 10362
rect 4551 10310 4603 10362
rect 4615 10310 4667 10362
rect 4679 10310 4731 10362
rect 11369 10310 11421 10362
rect 11433 10310 11485 10362
rect 11497 10310 11549 10362
rect 11561 10310 11613 10362
rect 11625 10310 11677 10362
rect 18315 10310 18367 10362
rect 18379 10310 18431 10362
rect 18443 10310 18495 10362
rect 18507 10310 18559 10362
rect 18571 10310 18623 10362
rect 25261 10310 25313 10362
rect 25325 10310 25377 10362
rect 25389 10310 25441 10362
rect 25453 10310 25505 10362
rect 25517 10310 25569 10362
rect 1584 10047 1636 10056
rect 1584 10013 1593 10047
rect 1593 10013 1627 10047
rect 1627 10013 1636 10047
rect 1584 10004 1636 10013
rect 7896 9766 7948 9818
rect 7960 9766 8012 9818
rect 8024 9766 8076 9818
rect 8088 9766 8140 9818
rect 8152 9766 8204 9818
rect 14842 9766 14894 9818
rect 14906 9766 14958 9818
rect 14970 9766 15022 9818
rect 15034 9766 15086 9818
rect 15098 9766 15150 9818
rect 21788 9766 21840 9818
rect 21852 9766 21904 9818
rect 21916 9766 21968 9818
rect 21980 9766 22032 9818
rect 22044 9766 22096 9818
rect 28734 9766 28786 9818
rect 28798 9766 28850 9818
rect 28862 9766 28914 9818
rect 28926 9766 28978 9818
rect 28990 9766 29042 9818
rect 28356 9435 28408 9444
rect 28356 9401 28365 9435
rect 28365 9401 28399 9435
rect 28399 9401 28408 9435
rect 28356 9392 28408 9401
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 4423 9222 4475 9274
rect 4487 9222 4539 9274
rect 4551 9222 4603 9274
rect 4615 9222 4667 9274
rect 4679 9222 4731 9274
rect 11369 9222 11421 9274
rect 11433 9222 11485 9274
rect 11497 9222 11549 9274
rect 11561 9222 11613 9274
rect 11625 9222 11677 9274
rect 18315 9222 18367 9274
rect 18379 9222 18431 9274
rect 18443 9222 18495 9274
rect 18507 9222 18559 9274
rect 18571 9222 18623 9274
rect 25261 9222 25313 9274
rect 25325 9222 25377 9274
rect 25389 9222 25441 9274
rect 25453 9222 25505 9274
rect 25517 9222 25569 9274
rect 28356 9095 28408 9104
rect 28356 9061 28365 9095
rect 28365 9061 28399 9095
rect 28399 9061 28408 9095
rect 28356 9052 28408 9061
rect 7896 8678 7948 8730
rect 7960 8678 8012 8730
rect 8024 8678 8076 8730
rect 8088 8678 8140 8730
rect 8152 8678 8204 8730
rect 14842 8678 14894 8730
rect 14906 8678 14958 8730
rect 14970 8678 15022 8730
rect 15034 8678 15086 8730
rect 15098 8678 15150 8730
rect 21788 8678 21840 8730
rect 21852 8678 21904 8730
rect 21916 8678 21968 8730
rect 21980 8678 22032 8730
rect 22044 8678 22096 8730
rect 28734 8678 28786 8730
rect 28798 8678 28850 8730
rect 28862 8678 28914 8730
rect 28926 8678 28978 8730
rect 28990 8678 29042 8730
rect 4423 8134 4475 8186
rect 4487 8134 4539 8186
rect 4551 8134 4603 8186
rect 4615 8134 4667 8186
rect 4679 8134 4731 8186
rect 11369 8134 11421 8186
rect 11433 8134 11485 8186
rect 11497 8134 11549 8186
rect 11561 8134 11613 8186
rect 11625 8134 11677 8186
rect 18315 8134 18367 8186
rect 18379 8134 18431 8186
rect 18443 8134 18495 8186
rect 18507 8134 18559 8186
rect 18571 8134 18623 8186
rect 25261 8134 25313 8186
rect 25325 8134 25377 8186
rect 25389 8134 25441 8186
rect 25453 8134 25505 8186
rect 25517 8134 25569 8186
rect 1584 7871 1636 7880
rect 1584 7837 1593 7871
rect 1593 7837 1627 7871
rect 1627 7837 1636 7871
rect 1584 7828 1636 7837
rect 28356 7871 28408 7880
rect 28356 7837 28365 7871
rect 28365 7837 28399 7871
rect 28399 7837 28408 7871
rect 28356 7828 28408 7837
rect 7896 7590 7948 7642
rect 7960 7590 8012 7642
rect 8024 7590 8076 7642
rect 8088 7590 8140 7642
rect 8152 7590 8204 7642
rect 14842 7590 14894 7642
rect 14906 7590 14958 7642
rect 14970 7590 15022 7642
rect 15034 7590 15086 7642
rect 15098 7590 15150 7642
rect 21788 7590 21840 7642
rect 21852 7590 21904 7642
rect 21916 7590 21968 7642
rect 21980 7590 22032 7642
rect 22044 7590 22096 7642
rect 28734 7590 28786 7642
rect 28798 7590 28850 7642
rect 28862 7590 28914 7642
rect 28926 7590 28978 7642
rect 28990 7590 29042 7642
rect 1584 7191 1636 7200
rect 1584 7157 1593 7191
rect 1593 7157 1627 7191
rect 1627 7157 1636 7191
rect 1584 7148 1636 7157
rect 4423 7046 4475 7098
rect 4487 7046 4539 7098
rect 4551 7046 4603 7098
rect 4615 7046 4667 7098
rect 4679 7046 4731 7098
rect 11369 7046 11421 7098
rect 11433 7046 11485 7098
rect 11497 7046 11549 7098
rect 11561 7046 11613 7098
rect 11625 7046 11677 7098
rect 18315 7046 18367 7098
rect 18379 7046 18431 7098
rect 18443 7046 18495 7098
rect 18507 7046 18559 7098
rect 18571 7046 18623 7098
rect 25261 7046 25313 7098
rect 25325 7046 25377 7098
rect 25389 7046 25441 7098
rect 25453 7046 25505 7098
rect 25517 7046 25569 7098
rect 28356 6783 28408 6792
rect 28356 6749 28365 6783
rect 28365 6749 28399 6783
rect 28399 6749 28408 6783
rect 28356 6740 28408 6749
rect 7896 6502 7948 6554
rect 7960 6502 8012 6554
rect 8024 6502 8076 6554
rect 8088 6502 8140 6554
rect 8152 6502 8204 6554
rect 14842 6502 14894 6554
rect 14906 6502 14958 6554
rect 14970 6502 15022 6554
rect 15034 6502 15086 6554
rect 15098 6502 15150 6554
rect 21788 6502 21840 6554
rect 21852 6502 21904 6554
rect 21916 6502 21968 6554
rect 21980 6502 22032 6554
rect 22044 6502 22096 6554
rect 28734 6502 28786 6554
rect 28798 6502 28850 6554
rect 28862 6502 28914 6554
rect 28926 6502 28978 6554
rect 28990 6502 29042 6554
rect 1584 6103 1636 6112
rect 1584 6069 1593 6103
rect 1593 6069 1627 6103
rect 1627 6069 1636 6103
rect 1584 6060 1636 6069
rect 4423 5958 4475 6010
rect 4487 5958 4539 6010
rect 4551 5958 4603 6010
rect 4615 5958 4667 6010
rect 4679 5958 4731 6010
rect 11369 5958 11421 6010
rect 11433 5958 11485 6010
rect 11497 5958 11549 6010
rect 11561 5958 11613 6010
rect 11625 5958 11677 6010
rect 18315 5958 18367 6010
rect 18379 5958 18431 6010
rect 18443 5958 18495 6010
rect 18507 5958 18559 6010
rect 18571 5958 18623 6010
rect 25261 5958 25313 6010
rect 25325 5958 25377 6010
rect 25389 5958 25441 6010
rect 25453 5958 25505 6010
rect 25517 5958 25569 6010
rect 28356 5695 28408 5704
rect 28356 5661 28365 5695
rect 28365 5661 28399 5695
rect 28399 5661 28408 5695
rect 28356 5652 28408 5661
rect 7896 5414 7948 5466
rect 7960 5414 8012 5466
rect 8024 5414 8076 5466
rect 8088 5414 8140 5466
rect 8152 5414 8204 5466
rect 14842 5414 14894 5466
rect 14906 5414 14958 5466
rect 14970 5414 15022 5466
rect 15034 5414 15086 5466
rect 15098 5414 15150 5466
rect 21788 5414 21840 5466
rect 21852 5414 21904 5466
rect 21916 5414 21968 5466
rect 21980 5414 22032 5466
rect 22044 5414 22096 5466
rect 28734 5414 28786 5466
rect 28798 5414 28850 5466
rect 28862 5414 28914 5466
rect 28926 5414 28978 5466
rect 28990 5414 29042 5466
rect 1584 5151 1636 5160
rect 1584 5117 1593 5151
rect 1593 5117 1627 5151
rect 1627 5117 1636 5151
rect 1584 5108 1636 5117
rect 28356 5015 28408 5024
rect 28356 4981 28365 5015
rect 28365 4981 28399 5015
rect 28399 4981 28408 5015
rect 28356 4972 28408 4981
rect 4423 4870 4475 4922
rect 4487 4870 4539 4922
rect 4551 4870 4603 4922
rect 4615 4870 4667 4922
rect 4679 4870 4731 4922
rect 11369 4870 11421 4922
rect 11433 4870 11485 4922
rect 11497 4870 11549 4922
rect 11561 4870 11613 4922
rect 11625 4870 11677 4922
rect 18315 4870 18367 4922
rect 18379 4870 18431 4922
rect 18443 4870 18495 4922
rect 18507 4870 18559 4922
rect 18571 4870 18623 4922
rect 25261 4870 25313 4922
rect 25325 4870 25377 4922
rect 25389 4870 25441 4922
rect 25453 4870 25505 4922
rect 25517 4870 25569 4922
rect 28356 4471 28408 4480
rect 28356 4437 28365 4471
rect 28365 4437 28399 4471
rect 28399 4437 28408 4471
rect 28356 4428 28408 4437
rect 7896 4326 7948 4378
rect 7960 4326 8012 4378
rect 8024 4326 8076 4378
rect 8088 4326 8140 4378
rect 8152 4326 8204 4378
rect 14842 4326 14894 4378
rect 14906 4326 14958 4378
rect 14970 4326 15022 4378
rect 15034 4326 15086 4378
rect 15098 4326 15150 4378
rect 21788 4326 21840 4378
rect 21852 4326 21904 4378
rect 21916 4326 21968 4378
rect 21980 4326 22032 4378
rect 22044 4326 22096 4378
rect 28734 4326 28786 4378
rect 28798 4326 28850 4378
rect 28862 4326 28914 4378
rect 28926 4326 28978 4378
rect 28990 4326 29042 4378
rect 17132 4020 17184 4072
rect 28356 4063 28408 4072
rect 28356 4029 28365 4063
rect 28365 4029 28399 4063
rect 28399 4029 28408 4063
rect 28356 4020 28408 4029
rect 1584 3927 1636 3936
rect 1584 3893 1593 3927
rect 1593 3893 1627 3927
rect 1627 3893 1636 3927
rect 1584 3884 1636 3893
rect 4423 3782 4475 3834
rect 4487 3782 4539 3834
rect 4551 3782 4603 3834
rect 4615 3782 4667 3834
rect 4679 3782 4731 3834
rect 11369 3782 11421 3834
rect 11433 3782 11485 3834
rect 11497 3782 11549 3834
rect 11561 3782 11613 3834
rect 11625 3782 11677 3834
rect 18315 3782 18367 3834
rect 18379 3782 18431 3834
rect 18443 3782 18495 3834
rect 18507 3782 18559 3834
rect 18571 3782 18623 3834
rect 25261 3782 25313 3834
rect 25325 3782 25377 3834
rect 25389 3782 25441 3834
rect 25453 3782 25505 3834
rect 25517 3782 25569 3834
rect 28356 3655 28408 3664
rect 28356 3621 28365 3655
rect 28365 3621 28399 3655
rect 28399 3621 28408 3655
rect 28356 3612 28408 3621
rect 1584 3519 1636 3528
rect 1584 3485 1593 3519
rect 1593 3485 1627 3519
rect 1627 3485 1636 3519
rect 1584 3476 1636 3485
rect 7896 3238 7948 3290
rect 7960 3238 8012 3290
rect 8024 3238 8076 3290
rect 8088 3238 8140 3290
rect 8152 3238 8204 3290
rect 14842 3238 14894 3290
rect 14906 3238 14958 3290
rect 14970 3238 15022 3290
rect 15034 3238 15086 3290
rect 15098 3238 15150 3290
rect 21788 3238 21840 3290
rect 21852 3238 21904 3290
rect 21916 3238 21968 3290
rect 21980 3238 22032 3290
rect 22044 3238 22096 3290
rect 28734 3238 28786 3290
rect 28798 3238 28850 3290
rect 28862 3238 28914 3290
rect 28926 3238 28978 3290
rect 28990 3238 29042 3290
rect 28356 2839 28408 2848
rect 28356 2805 28365 2839
rect 28365 2805 28399 2839
rect 28399 2805 28408 2839
rect 28356 2796 28408 2805
rect 4423 2694 4475 2746
rect 4487 2694 4539 2746
rect 4551 2694 4603 2746
rect 4615 2694 4667 2746
rect 4679 2694 4731 2746
rect 11369 2694 11421 2746
rect 11433 2694 11485 2746
rect 11497 2694 11549 2746
rect 11561 2694 11613 2746
rect 11625 2694 11677 2746
rect 18315 2694 18367 2746
rect 18379 2694 18431 2746
rect 18443 2694 18495 2746
rect 18507 2694 18559 2746
rect 18571 2694 18623 2746
rect 25261 2694 25313 2746
rect 25325 2694 25377 2746
rect 25389 2694 25441 2746
rect 25453 2694 25505 2746
rect 25517 2694 25569 2746
rect 7896 2150 7948 2202
rect 7960 2150 8012 2202
rect 8024 2150 8076 2202
rect 8088 2150 8140 2202
rect 8152 2150 8204 2202
rect 14842 2150 14894 2202
rect 14906 2150 14958 2202
rect 14970 2150 15022 2202
rect 15034 2150 15086 2202
rect 15098 2150 15150 2202
rect 21788 2150 21840 2202
rect 21852 2150 21904 2202
rect 21916 2150 21968 2202
rect 21980 2150 22032 2202
rect 22044 2150 22096 2202
rect 28734 2150 28786 2202
rect 28798 2150 28850 2202
rect 28862 2150 28914 2202
rect 28926 2150 28978 2202
rect 28990 2150 29042 2202
<< metal2 >>
rect 32 33238 520 33266
rect 32 25838 60 33238
rect 492 33130 520 33238
rect 570 33200 626 34000
rect 1674 33200 1730 34000
rect 2778 33200 2834 34000
rect 3882 33200 3938 34000
rect 4986 33200 5042 34000
rect 6090 33200 6146 34000
rect 6932 33238 7144 33266
rect 584 33130 612 33200
rect 492 33102 612 33130
rect 1688 28370 1716 33200
rect 2044 31272 2096 31278
rect 2044 31214 2096 31220
rect 2056 30734 2084 31214
rect 3056 31136 3108 31142
rect 3056 31078 3108 31084
rect 2044 30728 2096 30734
rect 2044 30670 2096 30676
rect 2688 30728 2740 30734
rect 2688 30670 2740 30676
rect 2044 30252 2096 30258
rect 2044 30194 2096 30200
rect 1952 29504 2004 29510
rect 1952 29446 2004 29452
rect 1964 29170 1992 29446
rect 1952 29164 2004 29170
rect 1952 29106 2004 29112
rect 1688 28342 1808 28370
rect 1674 28248 1730 28257
rect 1674 28183 1730 28192
rect 1584 26376 1636 26382
rect 1584 26318 1636 26324
rect 1596 26217 1624 26318
rect 1582 26208 1638 26217
rect 1582 26143 1638 26152
rect 1688 26042 1716 28183
rect 1780 26858 1808 28342
rect 2056 27985 2084 30194
rect 2700 30190 2728 30670
rect 3068 30326 3096 31078
rect 3056 30320 3108 30326
rect 2870 30288 2926 30297
rect 3056 30262 3108 30268
rect 3332 30252 3384 30258
rect 2870 30223 2926 30232
rect 2688 30184 2740 30190
rect 2318 30152 2374 30161
rect 2688 30126 2740 30132
rect 2318 30087 2374 30096
rect 2332 29306 2360 30087
rect 2700 29646 2728 30126
rect 2688 29640 2740 29646
rect 2594 29608 2650 29617
rect 2688 29582 2740 29588
rect 2594 29543 2596 29552
rect 2648 29543 2650 29552
rect 2596 29514 2648 29520
rect 2320 29300 2372 29306
rect 2320 29242 2372 29248
rect 2700 29238 2728 29582
rect 2688 29232 2740 29238
rect 2688 29174 2740 29180
rect 2136 29164 2188 29170
rect 2136 29106 2188 29112
rect 2042 27976 2098 27985
rect 2042 27911 2098 27920
rect 1768 26852 1820 26858
rect 1768 26794 1820 26800
rect 1676 26036 1728 26042
rect 1676 25978 1728 25984
rect 20 25832 72 25838
rect 20 25774 72 25780
rect 2148 25770 2176 29106
rect 2228 28960 2280 28966
rect 2228 28902 2280 28908
rect 2240 27441 2268 28902
rect 2700 28558 2728 29174
rect 2688 28552 2740 28558
rect 2688 28494 2740 28500
rect 2320 27872 2372 27878
rect 2320 27814 2372 27820
rect 2226 27432 2282 27441
rect 2226 27367 2282 27376
rect 2136 25764 2188 25770
rect 2136 25706 2188 25712
rect 2240 24954 2268 27367
rect 2332 26246 2360 27814
rect 2778 27568 2834 27577
rect 2596 27532 2648 27538
rect 2778 27503 2834 27512
rect 2596 27474 2648 27480
rect 2608 26450 2636 27474
rect 2596 26444 2648 26450
rect 2596 26386 2648 26392
rect 2608 26353 2636 26386
rect 2594 26344 2650 26353
rect 2594 26279 2650 26288
rect 2688 26308 2740 26314
rect 2688 26250 2740 26256
rect 2320 26240 2372 26246
rect 2318 26208 2320 26217
rect 2372 26208 2374 26217
rect 2318 26143 2374 26152
rect 2320 25696 2372 25702
rect 2320 25638 2372 25644
rect 2332 25537 2360 25638
rect 2318 25528 2374 25537
rect 2318 25463 2374 25472
rect 2228 24948 2280 24954
rect 2228 24890 2280 24896
rect 2700 24750 2728 26250
rect 2792 25430 2820 27503
rect 2884 27130 2912 30223
rect 3160 30212 3332 30240
rect 3056 30048 3108 30054
rect 3056 29990 3108 29996
rect 2962 29472 3018 29481
rect 2962 29407 3018 29416
rect 2872 27124 2924 27130
rect 2872 27066 2924 27072
rect 2872 26988 2924 26994
rect 2872 26930 2924 26936
rect 2780 25424 2832 25430
rect 2780 25366 2832 25372
rect 2884 24750 2912 26930
rect 2976 25498 3004 29407
rect 3068 29170 3096 29990
rect 3056 29164 3108 29170
rect 3056 29106 3108 29112
rect 3160 29050 3188 30212
rect 3332 30194 3384 30200
rect 3700 29504 3752 29510
rect 3700 29446 3752 29452
rect 3424 29300 3476 29306
rect 3424 29242 3476 29248
rect 3068 29022 3188 29050
rect 3068 26994 3096 29022
rect 3238 28656 3294 28665
rect 3238 28591 3294 28600
rect 3252 27130 3280 28591
rect 3436 27606 3464 29242
rect 3608 27940 3660 27946
rect 3608 27882 3660 27888
rect 3424 27600 3476 27606
rect 3424 27542 3476 27548
rect 3332 27464 3384 27470
rect 3332 27406 3384 27412
rect 3240 27124 3292 27130
rect 3240 27066 3292 27072
rect 3238 27024 3294 27033
rect 3056 26988 3108 26994
rect 3238 26959 3294 26968
rect 3056 26930 3108 26936
rect 3252 26518 3280 26959
rect 3240 26512 3292 26518
rect 3240 26454 3292 26460
rect 3240 26376 3292 26382
rect 3240 26318 3292 26324
rect 3056 26308 3108 26314
rect 3056 26250 3108 26256
rect 2964 25492 3016 25498
rect 2964 25434 3016 25440
rect 3068 25226 3096 26250
rect 3252 25809 3280 26318
rect 3238 25800 3294 25809
rect 3238 25735 3294 25744
rect 3056 25220 3108 25226
rect 3056 25162 3108 25168
rect 3252 24818 3280 25735
rect 3344 24857 3372 27406
rect 3620 27402 3648 27882
rect 3608 27396 3660 27402
rect 3608 27338 3660 27344
rect 3424 26784 3476 26790
rect 3424 26726 3476 26732
rect 3436 25362 3464 26726
rect 3620 26246 3648 27338
rect 3712 26897 3740 29446
rect 3792 27396 3844 27402
rect 3792 27338 3844 27344
rect 3804 26994 3832 27338
rect 3792 26988 3844 26994
rect 3792 26930 3844 26936
rect 3698 26888 3754 26897
rect 3698 26823 3754 26832
rect 3792 26308 3844 26314
rect 3792 26250 3844 26256
rect 3608 26240 3660 26246
rect 3608 26182 3660 26188
rect 3804 26081 3832 26250
rect 3790 26072 3846 26081
rect 3790 26007 3846 26016
rect 3896 25906 3924 33200
rect 4160 31680 4212 31686
rect 4160 31622 4212 31628
rect 4172 31346 4200 31622
rect 4160 31340 4212 31346
rect 4160 31282 4212 31288
rect 3976 31136 4028 31142
rect 3976 31078 4028 31084
rect 3988 29782 4016 31078
rect 4423 31036 4731 31045
rect 4423 31034 4429 31036
rect 4485 31034 4509 31036
rect 4565 31034 4589 31036
rect 4645 31034 4669 31036
rect 4725 31034 4731 31036
rect 4485 30982 4487 31034
rect 4667 30982 4669 31034
rect 4423 30980 4429 30982
rect 4485 30980 4509 30982
rect 4565 30980 4589 30982
rect 4645 30980 4669 30982
rect 4725 30980 4731 30982
rect 4423 30971 4731 30980
rect 4712 30796 4764 30802
rect 4712 30738 4764 30744
rect 4068 30660 4120 30666
rect 4068 30602 4120 30608
rect 4252 30660 4304 30666
rect 4252 30602 4304 30608
rect 3976 29776 4028 29782
rect 3976 29718 4028 29724
rect 4080 29510 4108 30602
rect 4160 30320 4212 30326
rect 4160 30262 4212 30268
rect 4068 29504 4120 29510
rect 4068 29446 4120 29452
rect 3976 28960 4028 28966
rect 3976 28902 4028 28908
rect 3988 28665 4016 28902
rect 3974 28656 4030 28665
rect 3974 28591 4030 28600
rect 4080 28506 4108 29446
rect 4172 28665 4200 30262
rect 4158 28656 4214 28665
rect 4158 28591 4214 28600
rect 3988 28478 4108 28506
rect 3988 27146 4016 28478
rect 4068 28416 4120 28422
rect 4068 28358 4120 28364
rect 4080 27470 4108 28358
rect 4160 27872 4212 27878
rect 4160 27814 4212 27820
rect 4068 27464 4120 27470
rect 4068 27406 4120 27412
rect 3988 27118 4108 27146
rect 3976 26988 4028 26994
rect 3976 26930 4028 26936
rect 3884 25900 3936 25906
rect 3884 25842 3936 25848
rect 3424 25356 3476 25362
rect 3424 25298 3476 25304
rect 3330 24848 3386 24857
rect 3240 24812 3292 24818
rect 3330 24783 3386 24792
rect 3240 24754 3292 24760
rect 2688 24744 2740 24750
rect 2688 24686 2740 24692
rect 2872 24744 2924 24750
rect 2872 24686 2924 24692
rect 2884 24410 2912 24686
rect 2872 24404 2924 24410
rect 2872 24346 2924 24352
rect 3988 24342 4016 26930
rect 4080 25702 4108 27118
rect 4172 26994 4200 27814
rect 4160 26988 4212 26994
rect 4160 26930 4212 26936
rect 4160 26784 4212 26790
rect 4160 26726 4212 26732
rect 4172 25974 4200 26726
rect 4160 25968 4212 25974
rect 4160 25910 4212 25916
rect 4068 25696 4120 25702
rect 4068 25638 4120 25644
rect 4264 25265 4292 30602
rect 4724 30598 4752 30738
rect 4344 30592 4396 30598
rect 4344 30534 4396 30540
rect 4712 30592 4764 30598
rect 4712 30534 4764 30540
rect 4356 26382 4384 30534
rect 4423 29948 4731 29957
rect 4423 29946 4429 29948
rect 4485 29946 4509 29948
rect 4565 29946 4589 29948
rect 4645 29946 4669 29948
rect 4725 29946 4731 29948
rect 4485 29894 4487 29946
rect 4667 29894 4669 29946
rect 4423 29892 4429 29894
rect 4485 29892 4509 29894
rect 4565 29892 4589 29894
rect 4645 29892 4669 29894
rect 4725 29892 4731 29894
rect 4423 29883 4731 29892
rect 4804 29776 4856 29782
rect 4804 29718 4856 29724
rect 4423 28860 4731 28869
rect 4423 28858 4429 28860
rect 4485 28858 4509 28860
rect 4565 28858 4589 28860
rect 4645 28858 4669 28860
rect 4725 28858 4731 28860
rect 4485 28806 4487 28858
rect 4667 28806 4669 28858
rect 4423 28804 4429 28806
rect 4485 28804 4509 28806
rect 4565 28804 4589 28806
rect 4645 28804 4669 28806
rect 4725 28804 4731 28806
rect 4423 28795 4731 28804
rect 4436 28484 4488 28490
rect 4436 28426 4488 28432
rect 4448 28082 4476 28426
rect 4436 28076 4488 28082
rect 4436 28018 4488 28024
rect 4423 27772 4731 27781
rect 4423 27770 4429 27772
rect 4485 27770 4509 27772
rect 4565 27770 4589 27772
rect 4645 27770 4669 27772
rect 4725 27770 4731 27772
rect 4485 27718 4487 27770
rect 4667 27718 4669 27770
rect 4423 27716 4429 27718
rect 4485 27716 4509 27718
rect 4565 27716 4589 27718
rect 4645 27716 4669 27718
rect 4725 27716 4731 27718
rect 4423 27707 4731 27716
rect 4816 27520 4844 29718
rect 4896 28076 4948 28082
rect 4896 28018 4948 28024
rect 4908 27674 4936 28018
rect 4896 27668 4948 27674
rect 4896 27610 4948 27616
rect 4816 27492 4936 27520
rect 4620 27464 4672 27470
rect 4672 27424 4844 27452
rect 4620 27406 4672 27412
rect 4712 27328 4764 27334
rect 4712 27270 4764 27276
rect 4724 27169 4752 27270
rect 4710 27160 4766 27169
rect 4710 27095 4766 27104
rect 4423 26684 4731 26693
rect 4423 26682 4429 26684
rect 4485 26682 4509 26684
rect 4565 26682 4589 26684
rect 4645 26682 4669 26684
rect 4725 26682 4731 26684
rect 4485 26630 4487 26682
rect 4667 26630 4669 26682
rect 4423 26628 4429 26630
rect 4485 26628 4509 26630
rect 4565 26628 4589 26630
rect 4645 26628 4669 26630
rect 4725 26628 4731 26630
rect 4423 26619 4731 26628
rect 4436 26512 4488 26518
rect 4434 26480 4436 26489
rect 4488 26480 4490 26489
rect 4434 26415 4490 26424
rect 4344 26376 4396 26382
rect 4344 26318 4396 26324
rect 4423 25596 4731 25605
rect 4423 25594 4429 25596
rect 4485 25594 4509 25596
rect 4565 25594 4589 25596
rect 4645 25594 4669 25596
rect 4725 25594 4731 25596
rect 4485 25542 4487 25594
rect 4667 25542 4669 25594
rect 4423 25540 4429 25542
rect 4485 25540 4509 25542
rect 4565 25540 4589 25542
rect 4645 25540 4669 25542
rect 4725 25540 4731 25542
rect 4423 25531 4731 25540
rect 4250 25256 4306 25265
rect 4250 25191 4306 25200
rect 4252 25152 4304 25158
rect 4252 25094 4304 25100
rect 4264 24818 4292 25094
rect 4252 24812 4304 24818
rect 4252 24754 4304 24760
rect 4816 24682 4844 27424
rect 4908 26042 4936 27492
rect 5000 26586 5028 33200
rect 6552 31680 6604 31686
rect 6552 31622 6604 31628
rect 5356 31476 5408 31482
rect 5356 31418 5408 31424
rect 5080 30796 5132 30802
rect 5080 30738 5132 30744
rect 4988 26580 5040 26586
rect 4988 26522 5040 26528
rect 4896 26036 4948 26042
rect 4896 25978 4948 25984
rect 4804 24676 4856 24682
rect 4804 24618 4856 24624
rect 4423 24508 4731 24517
rect 4423 24506 4429 24508
rect 4485 24506 4509 24508
rect 4565 24506 4589 24508
rect 4645 24506 4669 24508
rect 4725 24506 4731 24508
rect 4485 24454 4487 24506
rect 4667 24454 4669 24506
rect 4423 24452 4429 24454
rect 4485 24452 4509 24454
rect 4565 24452 4589 24454
rect 4645 24452 4669 24454
rect 4725 24452 4731 24454
rect 4423 24443 4731 24452
rect 4908 24410 4936 25978
rect 4988 25764 5040 25770
rect 4988 25706 5040 25712
rect 5000 25498 5028 25706
rect 4988 25492 5040 25498
rect 4988 25434 5040 25440
rect 5092 24818 5120 30738
rect 5172 29640 5224 29646
rect 5172 29582 5224 29588
rect 5184 27606 5212 29582
rect 5368 29170 5396 31418
rect 5540 31408 5592 31414
rect 5446 31376 5502 31385
rect 5540 31350 5592 31356
rect 5446 31311 5448 31320
rect 5500 31311 5502 31320
rect 5448 31282 5500 31288
rect 5552 30394 5580 31350
rect 6564 31346 6592 31622
rect 6552 31340 6604 31346
rect 6552 31282 6604 31288
rect 6276 31272 6328 31278
rect 6276 31214 6328 31220
rect 6642 31240 6698 31249
rect 6184 30728 6236 30734
rect 6184 30670 6236 30676
rect 5540 30388 5592 30394
rect 5540 30330 5592 30336
rect 5448 29232 5500 29238
rect 5552 29220 5580 30330
rect 6092 30320 6144 30326
rect 6090 30288 6092 30297
rect 6144 30288 6146 30297
rect 5908 30252 5960 30258
rect 6090 30223 6146 30232
rect 5908 30194 5960 30200
rect 5724 29708 5776 29714
rect 5724 29650 5776 29656
rect 5500 29192 5580 29220
rect 5448 29174 5500 29180
rect 5264 29164 5316 29170
rect 5264 29106 5316 29112
rect 5356 29164 5408 29170
rect 5356 29106 5408 29112
rect 5172 27600 5224 27606
rect 5172 27542 5224 27548
rect 5184 24993 5212 27542
rect 5276 25945 5304 29106
rect 5552 28762 5580 29192
rect 5540 28756 5592 28762
rect 5540 28698 5592 28704
rect 5448 28484 5500 28490
rect 5448 28426 5500 28432
rect 5356 27600 5408 27606
rect 5356 27542 5408 27548
rect 5368 27062 5396 27542
rect 5356 27056 5408 27062
rect 5356 26998 5408 27004
rect 5262 25936 5318 25945
rect 5262 25871 5318 25880
rect 5460 25430 5488 28426
rect 5552 28150 5580 28698
rect 5632 28212 5684 28218
rect 5632 28154 5684 28160
rect 5540 28144 5592 28150
rect 5540 28086 5592 28092
rect 5552 27470 5580 28086
rect 5540 27464 5592 27470
rect 5540 27406 5592 27412
rect 5644 26518 5672 28154
rect 5736 28082 5764 29650
rect 5816 28552 5868 28558
rect 5816 28494 5868 28500
rect 5828 28218 5856 28494
rect 5816 28212 5868 28218
rect 5816 28154 5868 28160
rect 5724 28076 5776 28082
rect 5724 28018 5776 28024
rect 5724 27532 5776 27538
rect 5724 27474 5776 27480
rect 5736 26761 5764 27474
rect 5722 26752 5778 26761
rect 5722 26687 5778 26696
rect 5724 26580 5776 26586
rect 5724 26522 5776 26528
rect 5632 26512 5684 26518
rect 5632 26454 5684 26460
rect 5538 26344 5594 26353
rect 5538 26279 5594 26288
rect 5552 26058 5580 26279
rect 5736 26058 5764 26522
rect 5552 26030 5764 26058
rect 5552 25906 5580 26030
rect 5632 25968 5684 25974
rect 5828 25956 5856 28154
rect 5684 25928 5856 25956
rect 5632 25910 5684 25916
rect 5540 25900 5592 25906
rect 5540 25842 5592 25848
rect 5920 25430 5948 30194
rect 6092 29844 6144 29850
rect 6092 29786 6144 29792
rect 6000 29300 6052 29306
rect 6000 29242 6052 29248
rect 6012 29209 6040 29242
rect 5998 29200 6054 29209
rect 5998 29135 6054 29144
rect 6104 27878 6132 29786
rect 6196 29170 6224 30670
rect 6288 29578 6316 31214
rect 6642 31175 6698 31184
rect 6656 30734 6684 31175
rect 6736 31136 6788 31142
rect 6736 31078 6788 31084
rect 6644 30728 6696 30734
rect 6644 30670 6696 30676
rect 6748 30433 6776 31078
rect 6734 30424 6790 30433
rect 6734 30359 6790 30368
rect 6644 30320 6696 30326
rect 6696 30268 6776 30274
rect 6644 30262 6776 30268
rect 6368 30252 6420 30258
rect 6656 30246 6776 30262
rect 6420 30212 6500 30240
rect 6368 30194 6420 30200
rect 6368 30048 6420 30054
rect 6368 29990 6420 29996
rect 6276 29572 6328 29578
rect 6276 29514 6328 29520
rect 6184 29164 6236 29170
rect 6184 29106 6236 29112
rect 6288 29050 6316 29514
rect 6380 29102 6408 29990
rect 6472 29306 6500 30212
rect 6644 30184 6696 30190
rect 6644 30126 6696 30132
rect 6460 29300 6512 29306
rect 6460 29242 6512 29248
rect 6196 29022 6316 29050
rect 6368 29096 6420 29102
rect 6368 29038 6420 29044
rect 6092 27872 6144 27878
rect 6092 27814 6144 27820
rect 6104 27674 6132 27814
rect 6092 27668 6144 27674
rect 6092 27610 6144 27616
rect 6000 27464 6052 27470
rect 6000 27406 6052 27412
rect 6012 26994 6040 27406
rect 6000 26988 6052 26994
rect 6000 26930 6052 26936
rect 6092 26920 6144 26926
rect 6196 26908 6224 29022
rect 6656 28994 6684 30126
rect 6748 29782 6776 30246
rect 6828 30048 6880 30054
rect 6828 29990 6880 29996
rect 6840 29850 6868 29990
rect 6828 29844 6880 29850
rect 6828 29786 6880 29792
rect 6736 29776 6788 29782
rect 6736 29718 6788 29724
rect 6828 29708 6880 29714
rect 6828 29650 6880 29656
rect 6840 28994 6868 29650
rect 6564 28966 6684 28994
rect 6748 28966 6868 28994
rect 6460 28756 6512 28762
rect 6460 28698 6512 28704
rect 6472 28014 6500 28698
rect 6460 28008 6512 28014
rect 6460 27950 6512 27956
rect 6368 27872 6420 27878
rect 6368 27814 6420 27820
rect 6274 27160 6330 27169
rect 6274 27095 6330 27104
rect 6144 26880 6224 26908
rect 6092 26862 6144 26868
rect 6000 26852 6052 26858
rect 6000 26794 6052 26800
rect 6012 26382 6040 26794
rect 6104 26586 6132 26862
rect 6092 26580 6144 26586
rect 6092 26522 6144 26528
rect 6092 26444 6144 26450
rect 6092 26386 6144 26392
rect 6000 26376 6052 26382
rect 6000 26318 6052 26324
rect 6012 26217 6040 26318
rect 5998 26208 6054 26217
rect 5998 26143 6054 26152
rect 6104 25770 6132 26386
rect 6288 26382 6316 27095
rect 6380 26994 6408 27814
rect 6472 27441 6500 27950
rect 6458 27432 6514 27441
rect 6458 27367 6460 27376
rect 6512 27367 6514 27376
rect 6460 27338 6512 27344
rect 6368 26988 6420 26994
rect 6368 26930 6420 26936
rect 6366 26752 6422 26761
rect 6366 26687 6422 26696
rect 6184 26376 6236 26382
rect 6184 26318 6236 26324
rect 6276 26376 6328 26382
rect 6276 26318 6328 26324
rect 6196 25906 6224 26318
rect 6276 26240 6328 26246
rect 6276 26182 6328 26188
rect 6288 25906 6316 26182
rect 6184 25900 6236 25906
rect 6184 25842 6236 25848
rect 6276 25900 6328 25906
rect 6276 25842 6328 25848
rect 6196 25786 6224 25842
rect 6092 25764 6144 25770
rect 6196 25758 6316 25786
rect 6092 25706 6144 25712
rect 5448 25424 5500 25430
rect 5448 25366 5500 25372
rect 5908 25424 5960 25430
rect 5908 25366 5960 25372
rect 5170 24984 5226 24993
rect 5170 24919 5226 24928
rect 5080 24812 5132 24818
rect 5080 24754 5132 24760
rect 4896 24404 4948 24410
rect 4896 24346 4948 24352
rect 3976 24336 4028 24342
rect 3976 24278 4028 24284
rect 1584 24200 1636 24206
rect 1582 24168 1584 24177
rect 1636 24168 1638 24177
rect 1582 24103 1638 24112
rect 5092 23798 5120 24754
rect 5460 24274 5488 25366
rect 6184 25288 6236 25294
rect 6184 25230 6236 25236
rect 6196 24954 6224 25230
rect 6184 24948 6236 24954
rect 6184 24890 6236 24896
rect 6288 24614 6316 25758
rect 6276 24608 6328 24614
rect 6276 24550 6328 24556
rect 5448 24268 5500 24274
rect 5448 24210 5500 24216
rect 5460 23866 5488 24210
rect 6380 24206 6408 26687
rect 6472 25537 6500 27338
rect 6564 26738 6592 28966
rect 6644 27396 6696 27402
rect 6644 27338 6696 27344
rect 6656 27130 6684 27338
rect 6644 27124 6696 27130
rect 6644 27066 6696 27072
rect 6748 26858 6776 28966
rect 6828 28688 6880 28694
rect 6828 28630 6880 28636
rect 6736 26852 6788 26858
rect 6736 26794 6788 26800
rect 6564 26710 6776 26738
rect 6642 26616 6698 26625
rect 6552 26580 6604 26586
rect 6642 26551 6698 26560
rect 6552 26522 6604 26528
rect 6564 25974 6592 26522
rect 6656 26518 6684 26551
rect 6644 26512 6696 26518
rect 6644 26454 6696 26460
rect 6748 26314 6776 26710
rect 6736 26308 6788 26314
rect 6736 26250 6788 26256
rect 6552 25968 6604 25974
rect 6552 25910 6604 25916
rect 6458 25528 6514 25537
rect 6458 25463 6514 25472
rect 6748 25226 6776 26250
rect 6460 25220 6512 25226
rect 6460 25162 6512 25168
rect 6736 25220 6788 25226
rect 6736 25162 6788 25168
rect 6472 24750 6500 25162
rect 6840 24750 6868 28630
rect 6932 25838 6960 33238
rect 7116 33130 7144 33238
rect 7194 33200 7250 34000
rect 8298 33200 8354 34000
rect 9402 33200 9458 34000
rect 10506 33200 10562 34000
rect 10612 33238 10824 33266
rect 7208 33130 7236 33200
rect 7116 33102 7236 33130
rect 7104 31680 7156 31686
rect 7104 31622 7156 31628
rect 7012 30320 7064 30326
rect 7010 30288 7012 30297
rect 7064 30288 7066 30297
rect 7010 30223 7066 30232
rect 7012 29776 7064 29782
rect 7012 29718 7064 29724
rect 7024 25838 7052 29718
rect 7116 28937 7144 31622
rect 7896 31580 8204 31589
rect 7896 31578 7902 31580
rect 7958 31578 7982 31580
rect 8038 31578 8062 31580
rect 8118 31578 8142 31580
rect 8198 31578 8204 31580
rect 7958 31526 7960 31578
rect 8140 31526 8142 31578
rect 7896 31524 7902 31526
rect 7958 31524 7982 31526
rect 8038 31524 8062 31526
rect 8118 31524 8142 31526
rect 8198 31524 8204 31526
rect 7896 31515 8204 31524
rect 7196 30932 7248 30938
rect 7196 30874 7248 30880
rect 7208 30705 7236 30874
rect 7562 30832 7618 30841
rect 7562 30767 7618 30776
rect 7194 30696 7250 30705
rect 7576 30666 7604 30767
rect 7194 30631 7250 30640
rect 7564 30660 7616 30666
rect 7208 29782 7236 30631
rect 7564 30602 7616 30608
rect 7656 30660 7708 30666
rect 7656 30602 7708 30608
rect 7288 30592 7340 30598
rect 7340 30540 7512 30546
rect 7288 30534 7512 30540
rect 7300 30518 7512 30534
rect 7288 30252 7340 30258
rect 7288 30194 7340 30200
rect 7196 29776 7248 29782
rect 7196 29718 7248 29724
rect 7300 29714 7328 30194
rect 7288 29708 7340 29714
rect 7288 29650 7340 29656
rect 7380 29572 7432 29578
rect 7380 29514 7432 29520
rect 7288 29300 7340 29306
rect 7288 29242 7340 29248
rect 7102 28928 7158 28937
rect 7102 28863 7158 28872
rect 7116 28490 7144 28863
rect 7104 28484 7156 28490
rect 7104 28426 7156 28432
rect 7116 28234 7144 28426
rect 7116 28206 7236 28234
rect 7104 28076 7156 28082
rect 7104 28018 7156 28024
rect 6920 25832 6972 25838
rect 6920 25774 6972 25780
rect 7012 25832 7064 25838
rect 7012 25774 7064 25780
rect 7116 25362 7144 28018
rect 7208 28014 7236 28206
rect 7196 28008 7248 28014
rect 7196 27950 7248 27956
rect 7196 27056 7248 27062
rect 7196 26998 7248 27004
rect 7208 26586 7236 26998
rect 7300 26586 7328 29242
rect 7196 26580 7248 26586
rect 7196 26522 7248 26528
rect 7288 26580 7340 26586
rect 7288 26522 7340 26528
rect 7300 26246 7328 26522
rect 7288 26240 7340 26246
rect 7288 26182 7340 26188
rect 7194 26072 7250 26081
rect 7194 26007 7250 26016
rect 7208 25770 7236 26007
rect 7196 25764 7248 25770
rect 7196 25706 7248 25712
rect 7104 25356 7156 25362
rect 7104 25298 7156 25304
rect 7116 24886 7144 25298
rect 7104 24880 7156 24886
rect 7104 24822 7156 24828
rect 6920 24812 6972 24818
rect 6920 24754 6972 24760
rect 6460 24744 6512 24750
rect 6460 24686 6512 24692
rect 6828 24744 6880 24750
rect 6828 24686 6880 24692
rect 6368 24200 6420 24206
rect 6368 24142 6420 24148
rect 6472 24070 6500 24686
rect 6932 24274 6960 24754
rect 7116 24274 7144 24822
rect 6920 24268 6972 24274
rect 6920 24210 6972 24216
rect 7104 24268 7156 24274
rect 7104 24210 7156 24216
rect 6460 24064 6512 24070
rect 6460 24006 6512 24012
rect 5448 23860 5500 23866
rect 5448 23802 5500 23808
rect 5080 23792 5132 23798
rect 5080 23734 5132 23740
rect 6472 23526 6500 24006
rect 6932 23866 6960 24210
rect 7392 23866 7420 29514
rect 7484 28370 7512 30518
rect 7668 30190 7696 30602
rect 7896 30492 8204 30501
rect 7896 30490 7902 30492
rect 7958 30490 7982 30492
rect 8038 30490 8062 30492
rect 8118 30490 8142 30492
rect 8198 30490 8204 30492
rect 7958 30438 7960 30490
rect 8140 30438 8142 30490
rect 7896 30436 7902 30438
rect 7958 30436 7982 30438
rect 8038 30436 8062 30438
rect 8118 30436 8142 30438
rect 8198 30436 8204 30438
rect 7896 30427 8204 30436
rect 7656 30184 7708 30190
rect 7656 30126 7708 30132
rect 7668 29306 7696 30126
rect 7748 29504 7800 29510
rect 7748 29446 7800 29452
rect 7656 29300 7708 29306
rect 7656 29242 7708 29248
rect 7760 29170 7788 29446
rect 7896 29404 8204 29413
rect 7896 29402 7902 29404
rect 7958 29402 7982 29404
rect 8038 29402 8062 29404
rect 8118 29402 8142 29404
rect 8198 29402 8204 29404
rect 7958 29350 7960 29402
rect 8140 29350 8142 29402
rect 7896 29348 7902 29350
rect 7958 29348 7982 29350
rect 8038 29348 8062 29350
rect 8118 29348 8142 29350
rect 8198 29348 8204 29350
rect 7896 29339 8204 29348
rect 7748 29164 7800 29170
rect 7748 29106 7800 29112
rect 7564 29096 7616 29102
rect 7562 29064 7564 29073
rect 7616 29064 7618 29073
rect 8312 29034 8340 33200
rect 10520 33130 10548 33200
rect 10612 33130 10640 33238
rect 10520 33102 10640 33130
rect 10796 31754 10824 33238
rect 11610 33200 11666 34000
rect 11716 33238 11928 33266
rect 11624 33130 11652 33200
rect 11716 33130 11744 33238
rect 11624 33102 11744 33130
rect 9312 31748 9364 31754
rect 10796 31726 11192 31754
rect 9312 31690 9364 31696
rect 8576 31680 8628 31686
rect 8576 31622 8628 31628
rect 8392 31136 8444 31142
rect 8392 31078 8444 31084
rect 8404 30394 8432 31078
rect 8588 30938 8616 31622
rect 8576 30932 8628 30938
rect 8576 30874 8628 30880
rect 9324 30734 9352 31690
rect 9680 31340 9732 31346
rect 9680 31282 9732 31288
rect 10048 31340 10100 31346
rect 10048 31282 10100 31288
rect 9404 31272 9456 31278
rect 9404 31214 9456 31220
rect 9220 30728 9272 30734
rect 9220 30670 9272 30676
rect 9312 30728 9364 30734
rect 9312 30670 9364 30676
rect 8392 30388 8444 30394
rect 8392 30330 8444 30336
rect 9036 30252 9088 30258
rect 9036 30194 9088 30200
rect 8944 30048 8996 30054
rect 8944 29990 8996 29996
rect 8484 29640 8536 29646
rect 8484 29582 8536 29588
rect 8390 29064 8446 29073
rect 7562 28999 7618 29008
rect 7748 29028 7800 29034
rect 7748 28970 7800 28976
rect 8300 29028 8352 29034
rect 8390 28999 8392 29008
rect 8300 28970 8352 28976
rect 8444 28999 8446 29008
rect 8392 28970 8444 28976
rect 7564 28416 7616 28422
rect 7484 28364 7564 28370
rect 7484 28358 7616 28364
rect 7484 28342 7604 28358
rect 7484 27674 7512 28342
rect 7656 28076 7708 28082
rect 7656 28018 7708 28024
rect 7564 27940 7616 27946
rect 7564 27882 7616 27888
rect 7472 27668 7524 27674
rect 7472 27610 7524 27616
rect 7576 27402 7604 27882
rect 7564 27396 7616 27402
rect 7564 27338 7616 27344
rect 7472 26376 7524 26382
rect 7576 26364 7604 27338
rect 7668 26625 7696 28018
rect 7654 26616 7710 26625
rect 7654 26551 7710 26560
rect 7656 26376 7708 26382
rect 7576 26336 7656 26364
rect 7472 26318 7524 26324
rect 7656 26318 7708 26324
rect 7484 25498 7512 26318
rect 7562 25528 7618 25537
rect 7472 25492 7524 25498
rect 7562 25463 7618 25472
rect 7472 25434 7524 25440
rect 7470 25392 7526 25401
rect 7470 25327 7526 25336
rect 7484 25226 7512 25327
rect 7472 25220 7524 25226
rect 7472 25162 7524 25168
rect 7484 24070 7512 25162
rect 7576 25158 7604 25463
rect 7564 25152 7616 25158
rect 7564 25094 7616 25100
rect 7562 24984 7618 24993
rect 7562 24919 7618 24928
rect 7576 24886 7604 24919
rect 7564 24880 7616 24886
rect 7564 24822 7616 24828
rect 7564 24608 7616 24614
rect 7564 24550 7616 24556
rect 7576 24138 7604 24550
rect 7668 24138 7696 26318
rect 7760 24682 7788 28970
rect 7896 28316 8204 28325
rect 7896 28314 7902 28316
rect 7958 28314 7982 28316
rect 8038 28314 8062 28316
rect 8118 28314 8142 28316
rect 8198 28314 8204 28316
rect 7958 28262 7960 28314
rect 8140 28262 8142 28314
rect 7896 28260 7902 28262
rect 7958 28260 7982 28262
rect 8038 28260 8062 28262
rect 8118 28260 8142 28262
rect 8198 28260 8204 28262
rect 7896 28251 8204 28260
rect 8300 28212 8352 28218
rect 8300 28154 8352 28160
rect 7896 27228 8204 27237
rect 7896 27226 7902 27228
rect 7958 27226 7982 27228
rect 8038 27226 8062 27228
rect 8118 27226 8142 27228
rect 8198 27226 8204 27228
rect 7958 27174 7960 27226
rect 8140 27174 8142 27226
rect 7896 27172 7902 27174
rect 7958 27172 7982 27174
rect 8038 27172 8062 27174
rect 8118 27172 8142 27174
rect 8198 27172 8204 27174
rect 7896 27163 8204 27172
rect 7896 26140 8204 26149
rect 7896 26138 7902 26140
rect 7958 26138 7982 26140
rect 8038 26138 8062 26140
rect 8118 26138 8142 26140
rect 8198 26138 8204 26140
rect 7958 26086 7960 26138
rect 8140 26086 8142 26138
rect 7896 26084 7902 26086
rect 7958 26084 7982 26086
rect 8038 26084 8062 26086
rect 8118 26084 8142 26086
rect 8198 26084 8204 26086
rect 7896 26075 8204 26084
rect 7840 25764 7892 25770
rect 7840 25706 7892 25712
rect 7852 25401 7880 25706
rect 8116 25696 8168 25702
rect 8116 25638 8168 25644
rect 7838 25392 7894 25401
rect 8128 25362 8156 25638
rect 7838 25327 7894 25336
rect 8116 25356 8168 25362
rect 8116 25298 8168 25304
rect 7896 25052 8204 25061
rect 7896 25050 7902 25052
rect 7958 25050 7982 25052
rect 8038 25050 8062 25052
rect 8118 25050 8142 25052
rect 8198 25050 8204 25052
rect 7958 24998 7960 25050
rect 8140 24998 8142 25050
rect 7896 24996 7902 24998
rect 7958 24996 7982 24998
rect 8038 24996 8062 24998
rect 8118 24996 8142 24998
rect 8198 24996 8204 24998
rect 7896 24987 8204 24996
rect 8312 24886 8340 28154
rect 8496 28150 8524 29582
rect 8576 29504 8628 29510
rect 8576 29446 8628 29452
rect 8588 28694 8616 29446
rect 8852 29164 8904 29170
rect 8852 29106 8904 29112
rect 8576 28688 8628 28694
rect 8576 28630 8628 28636
rect 8666 28656 8722 28665
rect 8666 28591 8722 28600
rect 8680 28490 8708 28591
rect 8576 28484 8628 28490
rect 8576 28426 8628 28432
rect 8668 28484 8720 28490
rect 8668 28426 8720 28432
rect 8484 28144 8536 28150
rect 8484 28086 8536 28092
rect 8496 27470 8524 28086
rect 8588 27878 8616 28426
rect 8576 27872 8628 27878
rect 8576 27814 8628 27820
rect 8484 27464 8536 27470
rect 8484 27406 8536 27412
rect 8758 27432 8814 27441
rect 8392 27328 8444 27334
rect 8392 27270 8444 27276
rect 8404 27130 8432 27270
rect 8392 27124 8444 27130
rect 8392 27066 8444 27072
rect 8496 26994 8524 27406
rect 8758 27367 8814 27376
rect 8668 27328 8720 27334
rect 8668 27270 8720 27276
rect 8680 27146 8708 27270
rect 8588 27118 8708 27146
rect 8588 26994 8616 27118
rect 8484 26988 8536 26994
rect 8484 26930 8536 26936
rect 8576 26988 8628 26994
rect 8576 26930 8628 26936
rect 8392 26920 8444 26926
rect 8392 26862 8444 26868
rect 8404 26790 8432 26862
rect 8392 26784 8444 26790
rect 8392 26726 8444 26732
rect 8392 26512 8444 26518
rect 8390 26480 8392 26489
rect 8444 26480 8446 26489
rect 8390 26415 8446 26424
rect 8496 26042 8524 26930
rect 8772 26625 8800 27367
rect 8758 26616 8814 26625
rect 8758 26551 8814 26560
rect 8864 26450 8892 29106
rect 8956 29073 8984 29990
rect 8942 29064 8998 29073
rect 8942 28999 8998 29008
rect 9048 27033 9076 30194
rect 9232 27452 9260 30670
rect 9312 27464 9364 27470
rect 9232 27424 9312 27452
rect 9312 27406 9364 27412
rect 9034 27024 9090 27033
rect 8944 26988 8996 26994
rect 9034 26959 9090 26968
rect 8944 26930 8996 26936
rect 8956 26466 8984 26930
rect 9128 26920 9180 26926
rect 9128 26862 9180 26868
rect 9036 26852 9088 26858
rect 9036 26794 9088 26800
rect 9048 26586 9076 26794
rect 9036 26580 9088 26586
rect 9036 26522 9088 26528
rect 8668 26444 8720 26450
rect 8668 26386 8720 26392
rect 8852 26444 8904 26450
rect 8956 26438 9076 26466
rect 9140 26450 9168 26862
rect 8852 26386 8904 26392
rect 8576 26308 8628 26314
rect 8576 26250 8628 26256
rect 8484 26036 8536 26042
rect 8484 25978 8536 25984
rect 8392 25288 8444 25294
rect 8392 25230 8444 25236
rect 8208 24880 8260 24886
rect 8208 24822 8260 24828
rect 8300 24880 8352 24886
rect 8300 24822 8352 24828
rect 8220 24750 8248 24822
rect 8208 24744 8260 24750
rect 8208 24686 8260 24692
rect 7748 24676 7800 24682
rect 7748 24618 7800 24624
rect 8404 24410 8432 25230
rect 8484 24608 8536 24614
rect 8484 24550 8536 24556
rect 8392 24404 8444 24410
rect 8392 24346 8444 24352
rect 8496 24206 8524 24550
rect 8484 24200 8536 24206
rect 8484 24142 8536 24148
rect 7564 24132 7616 24138
rect 7564 24074 7616 24080
rect 7656 24132 7708 24138
rect 7656 24074 7708 24080
rect 7472 24064 7524 24070
rect 7472 24006 7524 24012
rect 7896 23964 8204 23973
rect 7896 23962 7902 23964
rect 7958 23962 7982 23964
rect 8038 23962 8062 23964
rect 8118 23962 8142 23964
rect 8198 23962 8204 23964
rect 7958 23910 7960 23962
rect 8140 23910 8142 23962
rect 7896 23908 7902 23910
rect 7958 23908 7982 23910
rect 8038 23908 8062 23910
rect 8118 23908 8142 23910
rect 8198 23908 8204 23910
rect 7896 23899 8204 23908
rect 6920 23860 6972 23866
rect 6920 23802 6972 23808
rect 7380 23860 7432 23866
rect 7380 23802 7432 23808
rect 6932 23662 6960 23802
rect 8588 23730 8616 26250
rect 8680 24721 8708 26386
rect 8864 25362 8892 26386
rect 8944 26308 8996 26314
rect 8944 26250 8996 26256
rect 8956 25498 8984 26250
rect 8944 25492 8996 25498
rect 8944 25434 8996 25440
rect 9048 25430 9076 26438
rect 9128 26444 9180 26450
rect 9128 26386 9180 26392
rect 9128 26240 9180 26246
rect 9128 26182 9180 26188
rect 9036 25424 9088 25430
rect 9036 25366 9088 25372
rect 8852 25356 8904 25362
rect 8852 25298 8904 25304
rect 9140 25158 9168 26182
rect 9324 25770 9352 27406
rect 9416 27334 9444 31214
rect 9692 30297 9720 31282
rect 9772 31272 9824 31278
rect 9772 31214 9824 31220
rect 9784 30938 9812 31214
rect 10060 31142 10088 31282
rect 10048 31136 10100 31142
rect 10048 31078 10100 31084
rect 11060 31136 11112 31142
rect 11060 31078 11112 31084
rect 9772 30932 9824 30938
rect 9772 30874 9824 30880
rect 10968 30728 11020 30734
rect 11072 30716 11100 31078
rect 11164 30818 11192 31726
rect 11336 31476 11388 31482
rect 11336 31418 11388 31424
rect 11348 31142 11376 31418
rect 11336 31136 11388 31142
rect 11336 31078 11388 31084
rect 11794 31104 11850 31113
rect 11369 31036 11677 31045
rect 11794 31039 11850 31048
rect 11369 31034 11375 31036
rect 11431 31034 11455 31036
rect 11511 31034 11535 31036
rect 11591 31034 11615 31036
rect 11671 31034 11677 31036
rect 11431 30982 11433 31034
rect 11613 30982 11615 31034
rect 11369 30980 11375 30982
rect 11431 30980 11455 30982
rect 11511 30980 11535 30982
rect 11591 30980 11615 30982
rect 11671 30980 11677 30982
rect 11369 30971 11677 30980
rect 11336 30864 11388 30870
rect 11164 30812 11336 30818
rect 11164 30806 11388 30812
rect 11164 30790 11376 30806
rect 11072 30688 11284 30716
rect 11808 30705 11836 31039
rect 10968 30670 11020 30676
rect 10600 30660 10652 30666
rect 10600 30602 10652 30608
rect 10324 30388 10376 30394
rect 10324 30330 10376 30336
rect 10416 30388 10468 30394
rect 10416 30330 10468 30336
rect 9678 30288 9734 30297
rect 9678 30223 9734 30232
rect 9496 30184 9548 30190
rect 9496 30126 9548 30132
rect 9508 29646 9536 30126
rect 9680 29844 9732 29850
rect 9680 29786 9732 29792
rect 9496 29640 9548 29646
rect 9496 29582 9548 29588
rect 9588 29164 9640 29170
rect 9588 29106 9640 29112
rect 9600 28762 9628 29106
rect 9588 28756 9640 28762
rect 9588 28698 9640 28704
rect 9496 28688 9548 28694
rect 9496 28630 9548 28636
rect 9404 27328 9456 27334
rect 9404 27270 9456 27276
rect 9508 26586 9536 28630
rect 9600 28558 9628 28698
rect 9588 28552 9640 28558
rect 9588 28494 9640 28500
rect 9496 26580 9548 26586
rect 9496 26522 9548 26528
rect 9312 25764 9364 25770
rect 9312 25706 9364 25712
rect 9128 25152 9180 25158
rect 9128 25094 9180 25100
rect 8666 24712 8722 24721
rect 8666 24647 8722 24656
rect 8668 24404 8720 24410
rect 8668 24346 8720 24352
rect 8680 24206 8708 24346
rect 8668 24200 8720 24206
rect 9140 24188 9168 25094
rect 9508 24614 9536 26522
rect 9600 25974 9628 28494
rect 9692 28121 9720 29786
rect 10232 29640 10284 29646
rect 10232 29582 10284 29588
rect 9772 29572 9824 29578
rect 9772 29514 9824 29520
rect 9784 29238 9812 29514
rect 10244 29345 10272 29582
rect 10230 29336 10286 29345
rect 10230 29271 10286 29280
rect 9772 29232 9824 29238
rect 9772 29174 9824 29180
rect 9864 29164 9916 29170
rect 9864 29106 9916 29112
rect 9876 28937 9904 29106
rect 10336 28966 10364 30330
rect 10324 28960 10376 28966
rect 9862 28928 9918 28937
rect 10324 28902 10376 28908
rect 9862 28863 9918 28872
rect 9864 28620 9916 28626
rect 9864 28562 9916 28568
rect 9772 28552 9824 28558
rect 9772 28494 9824 28500
rect 9678 28112 9734 28121
rect 9678 28047 9734 28056
rect 9784 27062 9812 28494
rect 9772 27056 9824 27062
rect 9772 26998 9824 27004
rect 9876 26772 9904 28562
rect 9954 28248 10010 28257
rect 9954 28183 10010 28192
rect 9968 28150 9996 28183
rect 9956 28144 10008 28150
rect 9956 28086 10008 28092
rect 10140 27464 10192 27470
rect 10140 27406 10192 27412
rect 10152 27062 10180 27406
rect 10140 27056 10192 27062
rect 10140 26998 10192 27004
rect 9876 26744 9996 26772
rect 9680 26240 9732 26246
rect 9680 26182 9732 26188
rect 9588 25968 9640 25974
rect 9588 25910 9640 25916
rect 9692 25294 9720 26182
rect 9862 26072 9918 26081
rect 9862 26007 9918 26016
rect 9876 25906 9904 26007
rect 9864 25900 9916 25906
rect 9864 25842 9916 25848
rect 9864 25764 9916 25770
rect 9864 25706 9916 25712
rect 9770 25392 9826 25401
rect 9770 25327 9772 25336
rect 9824 25327 9826 25336
rect 9772 25298 9824 25304
rect 9876 25294 9904 25706
rect 9968 25294 9996 26744
rect 10048 26580 10100 26586
rect 10048 26522 10100 26528
rect 10060 25906 10088 26522
rect 10336 26450 10364 28902
rect 10324 26444 10376 26450
rect 10324 26386 10376 26392
rect 10322 26208 10378 26217
rect 10322 26143 10378 26152
rect 10336 25906 10364 26143
rect 10428 26081 10456 30330
rect 10508 29776 10560 29782
rect 10508 29718 10560 29724
rect 10414 26072 10470 26081
rect 10520 26042 10548 29718
rect 10612 26518 10640 30602
rect 10876 30592 10928 30598
rect 10876 30534 10928 30540
rect 10888 30376 10916 30534
rect 10980 30410 11008 30670
rect 11150 30560 11206 30569
rect 11150 30495 11206 30504
rect 10980 30382 11100 30410
rect 11164 30394 11192 30495
rect 10796 30348 10916 30376
rect 10692 30048 10744 30054
rect 10692 29990 10744 29996
rect 10704 29714 10732 29990
rect 10692 29708 10744 29714
rect 10692 29650 10744 29656
rect 10796 29594 10824 30348
rect 10876 30252 10928 30258
rect 10876 30194 10928 30200
rect 10704 29566 10824 29594
rect 10704 28422 10732 29566
rect 10784 29504 10836 29510
rect 10784 29446 10836 29452
rect 10692 28416 10744 28422
rect 10692 28358 10744 28364
rect 10704 26926 10732 28358
rect 10692 26920 10744 26926
rect 10692 26862 10744 26868
rect 10692 26784 10744 26790
rect 10796 26772 10824 29446
rect 10744 26744 10824 26772
rect 10692 26726 10744 26732
rect 10600 26512 10652 26518
rect 10600 26454 10652 26460
rect 10414 26007 10470 26016
rect 10508 26036 10560 26042
rect 10508 25978 10560 25984
rect 10048 25900 10100 25906
rect 10048 25842 10100 25848
rect 10324 25900 10376 25906
rect 10324 25842 10376 25848
rect 9680 25288 9732 25294
rect 9680 25230 9732 25236
rect 9864 25288 9916 25294
rect 9864 25230 9916 25236
rect 9956 25288 10008 25294
rect 9956 25230 10008 25236
rect 10598 25256 10654 25265
rect 9588 24880 9640 24886
rect 9692 24834 9720 25230
rect 9772 24948 9824 24954
rect 9772 24890 9824 24896
rect 9640 24828 9720 24834
rect 9588 24822 9720 24828
rect 9600 24806 9720 24822
rect 9588 24744 9640 24750
rect 9586 24712 9588 24721
rect 9640 24712 9642 24721
rect 9586 24647 9642 24656
rect 9496 24608 9548 24614
rect 9496 24550 9548 24556
rect 9600 24274 9628 24647
rect 9784 24410 9812 24890
rect 9772 24404 9824 24410
rect 9772 24346 9824 24352
rect 9588 24268 9640 24274
rect 9588 24210 9640 24216
rect 9220 24200 9272 24206
rect 9140 24160 9220 24188
rect 8668 24142 8720 24148
rect 9220 24142 9272 24148
rect 8576 23724 8628 23730
rect 8576 23666 8628 23672
rect 8680 23662 8708 24142
rect 6920 23656 6972 23662
rect 6920 23598 6972 23604
rect 8668 23656 8720 23662
rect 8668 23598 8720 23604
rect 1584 23520 1636 23526
rect 1582 23488 1584 23497
rect 6460 23520 6512 23526
rect 1636 23488 1638 23497
rect 6460 23462 6512 23468
rect 1582 23423 1638 23432
rect 4423 23420 4731 23429
rect 4423 23418 4429 23420
rect 4485 23418 4509 23420
rect 4565 23418 4589 23420
rect 4645 23418 4669 23420
rect 4725 23418 4731 23420
rect 4485 23366 4487 23418
rect 4667 23366 4669 23418
rect 4423 23364 4429 23366
rect 4485 23364 4509 23366
rect 4565 23364 4589 23366
rect 4645 23364 4669 23366
rect 4725 23364 4731 23366
rect 4423 23355 4731 23364
rect 9232 23322 9260 24142
rect 9600 23662 9628 24210
rect 9876 24206 9904 25230
rect 9968 24410 9996 25230
rect 10598 25191 10654 25200
rect 10612 25158 10640 25191
rect 10600 25152 10652 25158
rect 10600 25094 10652 25100
rect 10704 24818 10732 26726
rect 10416 24812 10468 24818
rect 10416 24754 10468 24760
rect 10692 24812 10744 24818
rect 10692 24754 10744 24760
rect 9956 24404 10008 24410
rect 9956 24346 10008 24352
rect 9864 24200 9916 24206
rect 9864 24142 9916 24148
rect 10428 24138 10456 24754
rect 10784 24608 10836 24614
rect 10784 24550 10836 24556
rect 10796 24206 10824 24550
rect 10888 24410 10916 30194
rect 11072 30190 11100 30382
rect 11152 30388 11204 30394
rect 11152 30330 11204 30336
rect 11060 30184 11112 30190
rect 11060 30126 11112 30132
rect 10968 30048 11020 30054
rect 10968 29990 11020 29996
rect 10980 29646 11008 29990
rect 10968 29640 11020 29646
rect 10968 29582 11020 29588
rect 11060 29232 11112 29238
rect 11060 29174 11112 29180
rect 11150 29200 11206 29209
rect 10968 29028 11020 29034
rect 10968 28970 11020 28976
rect 10980 28422 11008 28970
rect 10968 28416 11020 28422
rect 10968 28358 11020 28364
rect 10966 27568 11022 27577
rect 10966 27503 11022 27512
rect 10980 27470 11008 27503
rect 10968 27464 11020 27470
rect 10968 27406 11020 27412
rect 10968 26920 11020 26926
rect 10968 26862 11020 26868
rect 10980 26586 11008 26862
rect 10968 26580 11020 26586
rect 10968 26522 11020 26528
rect 10968 26444 11020 26450
rect 10968 26386 11020 26392
rect 10980 26246 11008 26386
rect 10968 26240 11020 26246
rect 10968 26182 11020 26188
rect 10980 26042 11008 26182
rect 10968 26036 11020 26042
rect 10968 25978 11020 25984
rect 10980 25430 11008 25978
rect 11072 25770 11100 29174
rect 11256 29170 11284 30688
rect 11794 30696 11850 30705
rect 11794 30631 11850 30640
rect 11794 30288 11850 30297
rect 11794 30223 11850 30232
rect 11704 30184 11756 30190
rect 11704 30126 11756 30132
rect 11369 29948 11677 29957
rect 11369 29946 11375 29948
rect 11431 29946 11455 29948
rect 11511 29946 11535 29948
rect 11591 29946 11615 29948
rect 11671 29946 11677 29948
rect 11431 29894 11433 29946
rect 11613 29894 11615 29946
rect 11369 29892 11375 29894
rect 11431 29892 11455 29894
rect 11511 29892 11535 29894
rect 11591 29892 11615 29894
rect 11671 29892 11677 29894
rect 11369 29883 11677 29892
rect 11716 29306 11744 30126
rect 11808 29782 11836 30223
rect 11796 29776 11848 29782
rect 11796 29718 11848 29724
rect 11704 29300 11756 29306
rect 11704 29242 11756 29248
rect 11150 29135 11206 29144
rect 11244 29164 11296 29170
rect 11164 25838 11192 29135
rect 11244 29106 11296 29112
rect 11336 29096 11388 29102
rect 11336 29038 11388 29044
rect 11348 28948 11376 29038
rect 11256 28920 11376 28948
rect 11256 26450 11284 28920
rect 11369 28860 11677 28869
rect 11369 28858 11375 28860
rect 11431 28858 11455 28860
rect 11511 28858 11535 28860
rect 11591 28858 11615 28860
rect 11671 28858 11677 28860
rect 11431 28806 11433 28858
rect 11613 28806 11615 28858
rect 11369 28804 11375 28806
rect 11431 28804 11455 28806
rect 11511 28804 11535 28806
rect 11591 28804 11615 28806
rect 11671 28804 11677 28806
rect 11369 28795 11677 28804
rect 11716 28014 11744 29242
rect 11808 29102 11836 29718
rect 11796 29096 11848 29102
rect 11796 29038 11848 29044
rect 11900 28966 11928 33238
rect 12714 33200 12770 34000
rect 13818 33200 13874 34000
rect 14922 33200 14978 34000
rect 16026 33200 16082 34000
rect 17130 33200 17186 34000
rect 18234 33200 18290 34000
rect 19338 33200 19394 34000
rect 20442 33200 20498 34000
rect 21546 33200 21602 34000
rect 22650 33200 22706 34000
rect 23754 33200 23810 34000
rect 24858 33200 24914 34000
rect 25962 33200 26018 34000
rect 27066 33200 27122 34000
rect 28170 33200 28226 34000
rect 29274 33200 29330 34000
rect 12532 31952 12584 31958
rect 12532 31894 12584 31900
rect 11980 31272 12032 31278
rect 11980 31214 12032 31220
rect 11992 29646 12020 31214
rect 12072 31204 12124 31210
rect 12072 31146 12124 31152
rect 12084 29753 12112 31146
rect 12164 30796 12216 30802
rect 12164 30738 12216 30744
rect 12176 30705 12204 30738
rect 12162 30696 12218 30705
rect 12162 30631 12218 30640
rect 12438 30016 12494 30025
rect 12438 29951 12494 29960
rect 12070 29744 12126 29753
rect 12070 29679 12126 29688
rect 11980 29640 12032 29646
rect 11980 29582 12032 29588
rect 11796 28960 11848 28966
rect 11796 28902 11848 28908
rect 11888 28960 11940 28966
rect 11888 28902 11940 28908
rect 11808 28801 11836 28902
rect 11794 28792 11850 28801
rect 11794 28727 11850 28736
rect 11794 28656 11850 28665
rect 11794 28591 11850 28600
rect 11704 28008 11756 28014
rect 11704 27950 11756 27956
rect 11369 27772 11677 27781
rect 11369 27770 11375 27772
rect 11431 27770 11455 27772
rect 11511 27770 11535 27772
rect 11591 27770 11615 27772
rect 11671 27770 11677 27772
rect 11431 27718 11433 27770
rect 11613 27718 11615 27770
rect 11369 27716 11375 27718
rect 11431 27716 11455 27718
rect 11511 27716 11535 27718
rect 11591 27716 11615 27718
rect 11671 27716 11677 27718
rect 11369 27707 11677 27716
rect 11612 27600 11664 27606
rect 11612 27542 11664 27548
rect 11624 26772 11652 27542
rect 11716 27538 11744 27950
rect 11704 27532 11756 27538
rect 11704 27474 11756 27480
rect 11624 26744 11744 26772
rect 11369 26684 11677 26693
rect 11369 26682 11375 26684
rect 11431 26682 11455 26684
rect 11511 26682 11535 26684
rect 11591 26682 11615 26684
rect 11671 26682 11677 26684
rect 11431 26630 11433 26682
rect 11613 26630 11615 26682
rect 11369 26628 11375 26630
rect 11431 26628 11455 26630
rect 11511 26628 11535 26630
rect 11591 26628 11615 26630
rect 11671 26628 11677 26630
rect 11369 26619 11677 26628
rect 11244 26444 11296 26450
rect 11244 26386 11296 26392
rect 11336 26376 11388 26382
rect 11336 26318 11388 26324
rect 11348 26042 11376 26318
rect 11716 26314 11744 26744
rect 11704 26308 11756 26314
rect 11704 26250 11756 26256
rect 11336 26036 11388 26042
rect 11336 25978 11388 25984
rect 11704 25968 11756 25974
rect 11702 25936 11704 25945
rect 11756 25936 11758 25945
rect 11702 25871 11758 25880
rect 11152 25832 11204 25838
rect 11152 25774 11204 25780
rect 11060 25764 11112 25770
rect 11060 25706 11112 25712
rect 11369 25596 11677 25605
rect 11369 25594 11375 25596
rect 11431 25594 11455 25596
rect 11511 25594 11535 25596
rect 11591 25594 11615 25596
rect 11671 25594 11677 25596
rect 11431 25542 11433 25594
rect 11613 25542 11615 25594
rect 11369 25540 11375 25542
rect 11431 25540 11455 25542
rect 11511 25540 11535 25542
rect 11591 25540 11615 25542
rect 11671 25540 11677 25542
rect 11369 25531 11677 25540
rect 10968 25424 11020 25430
rect 10968 25366 11020 25372
rect 11058 25392 11114 25401
rect 11058 25327 11114 25336
rect 11072 25294 11100 25327
rect 11808 25294 11836 28591
rect 11888 27600 11940 27606
rect 11888 27542 11940 27548
rect 11900 27402 11928 27542
rect 11888 27396 11940 27402
rect 11888 27338 11940 27344
rect 11060 25288 11112 25294
rect 11060 25230 11112 25236
rect 11152 25288 11204 25294
rect 11152 25230 11204 25236
rect 11796 25288 11848 25294
rect 11796 25230 11848 25236
rect 11164 24750 11192 25230
rect 11702 24848 11758 24857
rect 11702 24783 11758 24792
rect 11152 24744 11204 24750
rect 11152 24686 11204 24692
rect 10968 24676 11020 24682
rect 10968 24618 11020 24624
rect 10980 24410 11008 24618
rect 10876 24404 10928 24410
rect 10876 24346 10928 24352
rect 10968 24404 11020 24410
rect 10968 24346 11020 24352
rect 10784 24200 10836 24206
rect 10784 24142 10836 24148
rect 11164 24138 11192 24686
rect 11716 24682 11744 24783
rect 11704 24676 11756 24682
rect 11704 24618 11756 24624
rect 11369 24508 11677 24517
rect 11369 24506 11375 24508
rect 11431 24506 11455 24508
rect 11511 24506 11535 24508
rect 11591 24506 11615 24508
rect 11671 24506 11677 24508
rect 11431 24454 11433 24506
rect 11613 24454 11615 24506
rect 11369 24452 11375 24454
rect 11431 24452 11455 24454
rect 11511 24452 11535 24454
rect 11591 24452 11615 24454
rect 11671 24452 11677 24454
rect 11369 24443 11677 24452
rect 11808 24410 11836 25230
rect 11900 24818 11928 27338
rect 11992 26994 12020 29582
rect 12084 29238 12112 29679
rect 12164 29300 12216 29306
rect 12164 29242 12216 29248
rect 12256 29300 12308 29306
rect 12256 29242 12308 29248
rect 12072 29232 12124 29238
rect 12072 29174 12124 29180
rect 12176 28914 12204 29242
rect 12268 29034 12296 29242
rect 12348 29164 12400 29170
rect 12348 29106 12400 29112
rect 12256 29028 12308 29034
rect 12256 28970 12308 28976
rect 12084 28886 12204 28914
rect 12254 28928 12310 28937
rect 12084 28422 12112 28886
rect 12254 28863 12310 28872
rect 12268 28778 12296 28863
rect 12176 28750 12296 28778
rect 12360 28762 12388 29106
rect 12348 28756 12400 28762
rect 12176 28694 12204 28750
rect 12348 28698 12400 28704
rect 12164 28688 12216 28694
rect 12164 28630 12216 28636
rect 12256 28688 12308 28694
rect 12256 28630 12308 28636
rect 12268 28490 12296 28630
rect 12256 28484 12308 28490
rect 12256 28426 12308 28432
rect 12072 28416 12124 28422
rect 12072 28358 12124 28364
rect 12256 27668 12308 27674
rect 12256 27610 12308 27616
rect 12348 27668 12400 27674
rect 12348 27610 12400 27616
rect 12164 27464 12216 27470
rect 12164 27406 12216 27412
rect 11980 26988 12032 26994
rect 11980 26930 12032 26936
rect 12176 26042 12204 27406
rect 12268 27334 12296 27610
rect 12256 27328 12308 27334
rect 12256 27270 12308 27276
rect 12360 27010 12388 27610
rect 12452 27169 12480 29951
rect 12544 29306 12572 31894
rect 13832 31890 13860 33200
rect 14936 31958 14964 33200
rect 14924 31952 14976 31958
rect 14924 31894 14976 31900
rect 13820 31884 13872 31890
rect 13820 31826 13872 31832
rect 16120 31884 16172 31890
rect 16120 31826 16172 31832
rect 12992 31816 13044 31822
rect 12992 31758 13044 31764
rect 14554 31784 14610 31793
rect 13004 31346 13032 31758
rect 13636 31748 13688 31754
rect 13636 31690 13688 31696
rect 14280 31748 14332 31754
rect 14554 31719 14610 31728
rect 14280 31690 14332 31696
rect 13648 31482 13676 31690
rect 13636 31476 13688 31482
rect 13636 31418 13688 31424
rect 14096 31476 14148 31482
rect 14096 31418 14148 31424
rect 12992 31340 13044 31346
rect 12992 31282 13044 31288
rect 13084 31272 13136 31278
rect 13084 31214 13136 31220
rect 12714 30968 12770 30977
rect 12714 30903 12770 30912
rect 12992 30932 13044 30938
rect 12728 29578 12756 30903
rect 13096 30920 13124 31214
rect 13452 31136 13504 31142
rect 13452 31078 13504 31084
rect 13912 31136 13964 31142
rect 13912 31078 13964 31084
rect 13044 30892 13124 30920
rect 12992 30874 13044 30880
rect 12808 30388 12860 30394
rect 12808 30330 12860 30336
rect 12716 29572 12768 29578
rect 12716 29514 12768 29520
rect 12532 29300 12584 29306
rect 12532 29242 12584 29248
rect 12624 29232 12676 29238
rect 12624 29174 12676 29180
rect 12636 28490 12664 29174
rect 12716 28960 12768 28966
rect 12714 28928 12716 28937
rect 12768 28928 12770 28937
rect 12714 28863 12770 28872
rect 12624 28484 12676 28490
rect 12624 28426 12676 28432
rect 12636 27985 12664 28426
rect 12622 27976 12678 27985
rect 12622 27911 12678 27920
rect 12716 27940 12768 27946
rect 12716 27882 12768 27888
rect 12622 27840 12678 27849
rect 12622 27775 12678 27784
rect 12636 27470 12664 27775
rect 12624 27464 12676 27470
rect 12624 27406 12676 27412
rect 12728 27334 12756 27882
rect 12716 27328 12768 27334
rect 12716 27270 12768 27276
rect 12438 27160 12494 27169
rect 12438 27095 12494 27104
rect 12268 26982 12388 27010
rect 12164 26036 12216 26042
rect 12164 25978 12216 25984
rect 11978 25936 12034 25945
rect 11978 25871 12034 25880
rect 11992 25770 12020 25871
rect 11980 25764 12032 25770
rect 11980 25706 12032 25712
rect 12072 25696 12124 25702
rect 12072 25638 12124 25644
rect 12084 25498 12112 25638
rect 12072 25492 12124 25498
rect 12072 25434 12124 25440
rect 11980 25424 12032 25430
rect 11980 25366 12032 25372
rect 11992 25226 12020 25366
rect 11980 25220 12032 25226
rect 11980 25162 12032 25168
rect 11992 24818 12020 25162
rect 12072 25152 12124 25158
rect 12072 25094 12124 25100
rect 11888 24812 11940 24818
rect 11888 24754 11940 24760
rect 11980 24812 12032 24818
rect 11980 24754 12032 24760
rect 11796 24404 11848 24410
rect 11796 24346 11848 24352
rect 12084 24274 12112 25094
rect 12268 24614 12296 26982
rect 12440 26920 12492 26926
rect 12440 26862 12492 26868
rect 12348 26580 12400 26586
rect 12348 26522 12400 26528
rect 12360 26314 12388 26522
rect 12452 26466 12480 26862
rect 12532 26784 12584 26790
rect 12530 26752 12532 26761
rect 12584 26752 12586 26761
rect 12530 26687 12586 26696
rect 12544 26602 12572 26687
rect 12544 26574 12664 26602
rect 12728 26586 12756 27270
rect 12820 26926 12848 30330
rect 12900 30320 12952 30326
rect 12900 30262 12952 30268
rect 12912 29306 12940 30262
rect 13004 30258 13032 30874
rect 13360 30864 13412 30870
rect 13360 30806 13412 30812
rect 13268 30796 13320 30802
rect 13268 30738 13320 30744
rect 13280 30666 13308 30738
rect 13268 30660 13320 30666
rect 13268 30602 13320 30608
rect 12992 30252 13044 30258
rect 12992 30194 13044 30200
rect 13004 29696 13032 30194
rect 13084 30048 13136 30054
rect 13082 30016 13084 30025
rect 13136 30016 13138 30025
rect 13082 29951 13138 29960
rect 13174 29880 13230 29889
rect 13174 29815 13230 29824
rect 13084 29708 13136 29714
rect 13004 29668 13084 29696
rect 13084 29650 13136 29656
rect 12900 29300 12952 29306
rect 12900 29242 12952 29248
rect 13188 28994 13216 29815
rect 13268 29776 13320 29782
rect 13268 29718 13320 29724
rect 13096 28966 13216 28994
rect 12898 28928 12954 28937
rect 12898 28863 12954 28872
rect 12912 28218 12940 28863
rect 12900 28212 12952 28218
rect 12900 28154 12952 28160
rect 12992 28212 13044 28218
rect 12992 28154 13044 28160
rect 13004 27878 13032 28154
rect 12992 27872 13044 27878
rect 12992 27814 13044 27820
rect 13004 27418 13032 27814
rect 13096 27538 13124 28966
rect 13176 28620 13228 28626
rect 13176 28562 13228 28568
rect 13188 28529 13216 28562
rect 13174 28520 13230 28529
rect 13174 28455 13230 28464
rect 13176 28416 13228 28422
rect 13176 28358 13228 28364
rect 13188 28218 13216 28358
rect 13176 28212 13228 28218
rect 13176 28154 13228 28160
rect 13280 27962 13308 29718
rect 13372 28257 13400 30806
rect 13464 28762 13492 31078
rect 13636 30592 13688 30598
rect 13636 30534 13688 30540
rect 13648 30433 13676 30534
rect 13634 30424 13690 30433
rect 13634 30359 13690 30368
rect 13820 29844 13872 29850
rect 13820 29786 13872 29792
rect 13544 29504 13596 29510
rect 13544 29446 13596 29452
rect 13452 28756 13504 28762
rect 13452 28698 13504 28704
rect 13358 28248 13414 28257
rect 13358 28183 13414 28192
rect 13450 27976 13506 27985
rect 13280 27934 13400 27962
rect 13268 27872 13320 27878
rect 13268 27814 13320 27820
rect 13084 27532 13136 27538
rect 13084 27474 13136 27480
rect 13176 27464 13228 27470
rect 13174 27432 13176 27441
rect 13228 27432 13230 27441
rect 12900 27396 12952 27402
rect 13004 27390 13124 27418
rect 12900 27338 12952 27344
rect 12912 27130 12940 27338
rect 12992 27328 13044 27334
rect 12990 27296 12992 27305
rect 13044 27296 13046 27305
rect 12990 27231 13046 27240
rect 12990 27160 13046 27169
rect 12900 27124 12952 27130
rect 12990 27095 13046 27104
rect 12900 27066 12952 27072
rect 12808 26920 12860 26926
rect 12808 26862 12860 26868
rect 12452 26450 12572 26466
rect 12452 26444 12584 26450
rect 12452 26438 12532 26444
rect 12532 26386 12584 26392
rect 12440 26376 12492 26382
rect 12438 26344 12440 26353
rect 12492 26344 12494 26353
rect 12636 26330 12664 26574
rect 12716 26580 12768 26586
rect 12716 26522 12768 26528
rect 12348 26308 12400 26314
rect 12438 26279 12494 26288
rect 12544 26302 12664 26330
rect 12348 26250 12400 26256
rect 12544 25498 12572 26302
rect 13004 26194 13032 27095
rect 13096 26314 13124 27390
rect 13174 27367 13230 27376
rect 13174 27024 13230 27033
rect 13174 26959 13176 26968
rect 13228 26959 13230 26968
rect 13176 26930 13228 26936
rect 13084 26308 13136 26314
rect 13084 26250 13136 26256
rect 12912 26166 13032 26194
rect 13176 26240 13228 26246
rect 13176 26182 13228 26188
rect 12624 25968 12676 25974
rect 12676 25916 12756 25922
rect 12624 25910 12756 25916
rect 12636 25894 12756 25910
rect 12622 25800 12678 25809
rect 12622 25735 12678 25744
rect 12636 25702 12664 25735
rect 12728 25702 12756 25894
rect 12624 25696 12676 25702
rect 12624 25638 12676 25644
rect 12716 25696 12768 25702
rect 12716 25638 12768 25644
rect 12532 25492 12584 25498
rect 12532 25434 12584 25440
rect 12348 25220 12400 25226
rect 12636 25208 12664 25638
rect 12716 25220 12768 25226
rect 12636 25180 12716 25208
rect 12348 25162 12400 25168
rect 12716 25162 12768 25168
rect 12360 24954 12388 25162
rect 12348 24948 12400 24954
rect 12348 24890 12400 24896
rect 12912 24818 12940 26166
rect 12990 26072 13046 26081
rect 12990 26007 13046 26016
rect 13004 25974 13032 26007
rect 12992 25968 13044 25974
rect 12992 25910 13044 25916
rect 13188 25906 13216 26182
rect 13176 25900 13228 25906
rect 13176 25842 13228 25848
rect 13084 25832 13136 25838
rect 13084 25774 13136 25780
rect 13096 25294 13124 25774
rect 13280 25702 13308 27814
rect 13372 26314 13400 27934
rect 13450 27911 13506 27920
rect 13464 27878 13492 27911
rect 13452 27872 13504 27878
rect 13452 27814 13504 27820
rect 13452 27464 13504 27470
rect 13452 27406 13504 27412
rect 13464 27305 13492 27406
rect 13450 27296 13506 27305
rect 13450 27231 13506 27240
rect 13464 26897 13492 27231
rect 13556 27130 13584 29446
rect 13832 28994 13860 29786
rect 13924 29578 13952 31078
rect 14004 30796 14056 30802
rect 14004 30738 14056 30744
rect 13912 29572 13964 29578
rect 13912 29514 13964 29520
rect 13832 28966 13952 28994
rect 13636 28620 13688 28626
rect 13636 28562 13688 28568
rect 13544 27124 13596 27130
rect 13544 27066 13596 27072
rect 13648 27062 13676 28562
rect 13924 28529 13952 28966
rect 14016 28558 14044 30738
rect 14108 28762 14136 31418
rect 14188 31408 14240 31414
rect 14188 31350 14240 31356
rect 14200 30938 14228 31350
rect 14188 30932 14240 30938
rect 14188 30874 14240 30880
rect 14292 30705 14320 31690
rect 14568 31686 14596 31719
rect 14556 31680 14608 31686
rect 14556 31622 14608 31628
rect 14568 31414 14596 31622
rect 14842 31580 15150 31589
rect 14842 31578 14848 31580
rect 14904 31578 14928 31580
rect 14984 31578 15008 31580
rect 15064 31578 15088 31580
rect 15144 31578 15150 31580
rect 14904 31526 14906 31578
rect 15086 31526 15088 31578
rect 14842 31524 14848 31526
rect 14904 31524 14928 31526
rect 14984 31524 15008 31526
rect 15064 31524 15088 31526
rect 15144 31524 15150 31526
rect 14842 31515 15150 31524
rect 14556 31408 14608 31414
rect 14476 31368 14556 31396
rect 14278 30696 14334 30705
rect 14278 30631 14334 30640
rect 14188 30320 14240 30326
rect 14188 30262 14240 30268
rect 14200 29209 14228 30262
rect 14186 29200 14242 29209
rect 14186 29135 14242 29144
rect 14096 28756 14148 28762
rect 14096 28698 14148 28704
rect 14108 28665 14136 28698
rect 14094 28656 14150 28665
rect 14292 28626 14320 30631
rect 14372 30592 14424 30598
rect 14372 30534 14424 30540
rect 14384 30394 14412 30534
rect 14372 30388 14424 30394
rect 14372 30330 14424 30336
rect 14476 29782 14504 31368
rect 14556 31350 14608 31356
rect 16132 31346 16160 31826
rect 16396 31816 16448 31822
rect 16396 31758 16448 31764
rect 15660 31340 15712 31346
rect 15660 31282 15712 31288
rect 16120 31340 16172 31346
rect 16120 31282 16172 31288
rect 15568 31136 15620 31142
rect 15568 31078 15620 31084
rect 15382 30968 15438 30977
rect 15382 30903 15438 30912
rect 14556 30864 14608 30870
rect 14556 30806 14608 30812
rect 14568 30666 14596 30806
rect 15396 30734 15424 30903
rect 15108 30728 15160 30734
rect 15384 30728 15436 30734
rect 15160 30688 15332 30716
rect 15108 30670 15160 30676
rect 14556 30660 14608 30666
rect 14556 30602 14608 30608
rect 15304 30580 15332 30688
rect 15384 30670 15436 30676
rect 15304 30552 15424 30580
rect 14842 30492 15150 30501
rect 14842 30490 14848 30492
rect 14904 30490 14928 30492
rect 14984 30490 15008 30492
rect 15064 30490 15088 30492
rect 15144 30490 15150 30492
rect 14904 30438 14906 30490
rect 15086 30438 15088 30490
rect 14842 30436 14848 30438
rect 14904 30436 14928 30438
rect 14984 30436 15008 30438
rect 15064 30436 15088 30438
rect 15144 30436 15150 30438
rect 14554 30424 14610 30433
rect 14842 30427 15150 30436
rect 15396 30410 15424 30552
rect 15580 30433 15608 31078
rect 15672 30802 15700 31282
rect 16120 30864 16172 30870
rect 16120 30806 16172 30812
rect 15660 30796 15712 30802
rect 15660 30738 15712 30744
rect 15566 30424 15622 30433
rect 15396 30382 15433 30410
rect 14554 30359 14610 30368
rect 14568 30002 14596 30359
rect 14832 30320 14884 30326
rect 15405 30274 15433 30382
rect 15566 30359 15622 30368
rect 14832 30262 14884 30268
rect 14568 29974 14780 30002
rect 14464 29776 14516 29782
rect 14464 29718 14516 29724
rect 14568 29646 14596 29974
rect 14646 29880 14702 29889
rect 14752 29850 14780 29974
rect 14844 29889 14872 30262
rect 14924 30252 14976 30258
rect 14924 30194 14976 30200
rect 15396 30246 15433 30274
rect 15660 30320 15712 30326
rect 15660 30262 15712 30268
rect 15476 30252 15528 30258
rect 14830 29880 14886 29889
rect 14646 29815 14702 29824
rect 14740 29844 14792 29850
rect 14556 29640 14608 29646
rect 14660 29628 14688 29815
rect 14830 29815 14886 29824
rect 14740 29786 14792 29792
rect 14936 29714 14964 30194
rect 15108 30116 15160 30122
rect 15028 30076 15108 30104
rect 15028 29753 15056 30076
rect 15108 30058 15160 30064
rect 15200 30048 15252 30054
rect 15396 30036 15424 30246
rect 15476 30194 15528 30200
rect 15200 29990 15252 29996
rect 15304 30008 15424 30036
rect 15014 29744 15070 29753
rect 14924 29708 14976 29714
rect 15212 29714 15240 29990
rect 15304 29850 15332 30008
rect 15292 29844 15344 29850
rect 15292 29786 15344 29792
rect 15384 29844 15436 29850
rect 15488 29832 15516 30194
rect 15672 30122 15700 30262
rect 15660 30116 15712 30122
rect 15660 30058 15712 30064
rect 15764 29850 15976 29866
rect 15752 29844 15976 29850
rect 15488 29804 15608 29832
rect 15384 29786 15436 29792
rect 15405 29714 15433 29786
rect 15474 29744 15530 29753
rect 15014 29679 15070 29688
rect 15108 29708 15160 29714
rect 14924 29650 14976 29656
rect 15108 29650 15160 29656
rect 15200 29708 15252 29714
rect 15200 29650 15252 29656
rect 15292 29708 15344 29714
rect 15292 29650 15344 29656
rect 15384 29708 15436 29714
rect 15474 29679 15530 29688
rect 15384 29650 15436 29656
rect 14740 29640 14792 29646
rect 14660 29600 14740 29628
rect 14556 29582 14608 29588
rect 14740 29582 14792 29588
rect 15120 29594 15148 29650
rect 15120 29566 15240 29594
rect 15304 29578 15332 29650
rect 14648 29504 14700 29510
rect 14646 29472 14648 29481
rect 14700 29472 14702 29481
rect 14646 29407 14702 29416
rect 14842 29404 15150 29413
rect 14842 29402 14848 29404
rect 14904 29402 14928 29404
rect 14984 29402 15008 29404
rect 15064 29402 15088 29404
rect 15144 29402 15150 29404
rect 14904 29350 14906 29402
rect 15086 29350 15088 29402
rect 14842 29348 14848 29350
rect 14904 29348 14928 29350
rect 14984 29348 15008 29350
rect 15064 29348 15088 29350
rect 15144 29348 15150 29350
rect 14842 29339 15150 29348
rect 14464 29300 14516 29306
rect 14464 29242 14516 29248
rect 14832 29300 14884 29306
rect 14832 29242 14884 29248
rect 14094 28591 14150 28600
rect 14280 28620 14332 28626
rect 14280 28562 14332 28568
rect 14004 28552 14056 28558
rect 13910 28520 13966 28529
rect 13820 28484 13872 28490
rect 14004 28494 14056 28500
rect 13910 28455 13966 28464
rect 14096 28484 14148 28490
rect 13820 28426 13872 28432
rect 14096 28426 14148 28432
rect 13728 28416 13780 28422
rect 13728 28358 13780 28364
rect 13832 28370 13860 28426
rect 13636 27056 13688 27062
rect 13636 26998 13688 27004
rect 13450 26888 13506 26897
rect 13740 26874 13768 28358
rect 13832 28342 14044 28370
rect 13912 27872 13964 27878
rect 13912 27814 13964 27820
rect 13818 27704 13874 27713
rect 13818 27639 13874 27648
rect 13832 27538 13860 27639
rect 13820 27532 13872 27538
rect 13820 27474 13872 27480
rect 13924 27441 13952 27814
rect 13910 27432 13966 27441
rect 14016 27402 14044 28342
rect 13910 27367 13966 27376
rect 14004 27396 14056 27402
rect 14004 27338 14056 27344
rect 13820 27328 13872 27334
rect 13820 27270 13872 27276
rect 13450 26823 13506 26832
rect 13648 26846 13768 26874
rect 13648 26586 13676 26846
rect 13636 26580 13688 26586
rect 13636 26522 13688 26528
rect 13634 26480 13690 26489
rect 13452 26444 13504 26450
rect 13634 26415 13636 26424
rect 13452 26386 13504 26392
rect 13688 26415 13690 26424
rect 13636 26386 13688 26392
rect 13360 26308 13412 26314
rect 13360 26250 13412 26256
rect 13268 25696 13320 25702
rect 13268 25638 13320 25644
rect 13084 25288 13136 25294
rect 13084 25230 13136 25236
rect 13372 24818 13400 26250
rect 13464 25922 13492 26386
rect 13464 25906 13584 25922
rect 13464 25900 13596 25906
rect 13464 25894 13544 25900
rect 13544 25842 13596 25848
rect 13832 24886 13860 27270
rect 14016 27062 14044 27338
rect 14004 27056 14056 27062
rect 14108 27033 14136 28426
rect 14372 28008 14424 28014
rect 14372 27950 14424 27956
rect 14280 27872 14332 27878
rect 14280 27814 14332 27820
rect 14186 27704 14242 27713
rect 14186 27639 14242 27648
rect 14004 26998 14056 27004
rect 14094 27024 14150 27033
rect 13912 26512 13964 26518
rect 13912 26454 13964 26460
rect 13924 25906 13952 26454
rect 13912 25900 13964 25906
rect 13912 25842 13964 25848
rect 14016 25158 14044 26998
rect 14094 26959 14150 26968
rect 14108 26790 14136 26959
rect 14096 26784 14148 26790
rect 14096 26726 14148 26732
rect 14096 26580 14148 26586
rect 14096 26522 14148 26528
rect 14108 26353 14136 26522
rect 14200 26382 14228 27639
rect 14292 26858 14320 27814
rect 14384 27606 14412 27950
rect 14476 27606 14504 29242
rect 14844 29186 14872 29242
rect 14660 29158 14872 29186
rect 15108 29164 15160 29170
rect 14660 27606 14688 29158
rect 15212 29152 15240 29566
rect 15292 29572 15344 29578
rect 15292 29514 15344 29520
rect 15304 29238 15332 29514
rect 15382 29336 15438 29345
rect 15382 29271 15384 29280
rect 15436 29271 15438 29280
rect 15384 29242 15436 29248
rect 15292 29232 15344 29238
rect 15292 29174 15344 29180
rect 15160 29124 15240 29152
rect 15108 29106 15160 29112
rect 14924 29096 14976 29102
rect 14738 29064 14794 29073
rect 14924 29038 14976 29044
rect 14738 28999 14794 29008
rect 14752 28626 14780 28999
rect 14936 28626 14964 29038
rect 15028 29034 15240 29050
rect 15016 29028 15240 29034
rect 15068 29022 15240 29028
rect 15016 28970 15068 28976
rect 14740 28620 14792 28626
rect 14740 28562 14792 28568
rect 14924 28620 14976 28626
rect 14924 28562 14976 28568
rect 14842 28316 15150 28325
rect 14842 28314 14848 28316
rect 14904 28314 14928 28316
rect 14984 28314 15008 28316
rect 15064 28314 15088 28316
rect 15144 28314 15150 28316
rect 14904 28262 14906 28314
rect 15086 28262 15088 28314
rect 14842 28260 14848 28262
rect 14904 28260 14928 28262
rect 14984 28260 15008 28262
rect 15064 28260 15088 28262
rect 15144 28260 15150 28262
rect 14842 28251 15150 28260
rect 15014 28112 15070 28121
rect 14740 28076 14792 28082
rect 15014 28047 15016 28056
rect 14740 28018 14792 28024
rect 15068 28047 15070 28056
rect 15016 28018 15068 28024
rect 14372 27600 14424 27606
rect 14372 27542 14424 27548
rect 14464 27600 14516 27606
rect 14464 27542 14516 27548
rect 14648 27600 14700 27606
rect 14648 27542 14700 27548
rect 14384 27130 14412 27542
rect 14660 27452 14688 27542
rect 14476 27424 14688 27452
rect 14372 27124 14424 27130
rect 14372 27066 14424 27072
rect 14476 26994 14504 27424
rect 14464 26988 14516 26994
rect 14464 26930 14516 26936
rect 14752 26858 14780 28018
rect 15108 27940 15160 27946
rect 15108 27882 15160 27888
rect 15120 27674 15148 27882
rect 15108 27668 15160 27674
rect 15108 27610 15160 27616
rect 15108 27532 15160 27538
rect 15108 27474 15160 27480
rect 15120 27334 15148 27474
rect 15108 27328 15160 27334
rect 15108 27270 15160 27276
rect 14842 27228 15150 27237
rect 14842 27226 14848 27228
rect 14904 27226 14928 27228
rect 14984 27226 15008 27228
rect 15064 27226 15088 27228
rect 15144 27226 15150 27228
rect 14904 27174 14906 27226
rect 15086 27174 15088 27226
rect 14842 27172 14848 27174
rect 14904 27172 14928 27174
rect 14984 27172 15008 27174
rect 15064 27172 15088 27174
rect 15144 27172 15150 27174
rect 14842 27163 15150 27172
rect 15212 27130 15240 29022
rect 15304 27674 15332 29174
rect 15384 28960 15436 28966
rect 15384 28902 15436 28908
rect 15396 27878 15424 28902
rect 15488 28762 15516 29679
rect 15580 29560 15608 29804
rect 15804 29838 15976 29844
rect 15752 29786 15804 29792
rect 15948 29782 15976 29838
rect 15844 29776 15896 29782
rect 15844 29718 15896 29724
rect 15936 29776 15988 29782
rect 15936 29718 15988 29724
rect 15856 29617 15884 29718
rect 15548 29532 15608 29560
rect 15842 29608 15898 29617
rect 15842 29543 15898 29552
rect 16028 29572 16080 29578
rect 15548 29322 15576 29532
rect 16028 29514 16080 29520
rect 15548 29294 15700 29322
rect 15476 28756 15528 28762
rect 15476 28698 15528 28704
rect 15476 28008 15528 28014
rect 15474 27976 15476 27985
rect 15528 27976 15530 27985
rect 15474 27911 15530 27920
rect 15384 27872 15436 27878
rect 15384 27814 15436 27820
rect 15292 27668 15344 27674
rect 15292 27610 15344 27616
rect 15292 27328 15344 27334
rect 15292 27270 15344 27276
rect 15200 27124 15252 27130
rect 15200 27066 15252 27072
rect 14832 26988 14884 26994
rect 14832 26930 14884 26936
rect 14280 26852 14332 26858
rect 14280 26794 14332 26800
rect 14740 26852 14792 26858
rect 14740 26794 14792 26800
rect 14188 26376 14240 26382
rect 14094 26344 14150 26353
rect 14188 26318 14240 26324
rect 14094 26279 14150 26288
rect 14292 25430 14320 26794
rect 14462 26752 14518 26761
rect 14844 26738 14872 26930
rect 15304 26926 15332 27270
rect 15292 26920 15344 26926
rect 15292 26862 15344 26868
rect 14462 26687 14518 26696
rect 14752 26710 14872 26738
rect 14476 26382 14504 26687
rect 14464 26376 14516 26382
rect 14464 26318 14516 26324
rect 14476 26246 14504 26318
rect 14464 26240 14516 26246
rect 14464 26182 14516 26188
rect 14752 25974 14780 26710
rect 15304 26518 15332 26862
rect 15292 26512 15344 26518
rect 15292 26454 15344 26460
rect 14842 26140 15150 26149
rect 14842 26138 14848 26140
rect 14904 26138 14928 26140
rect 14984 26138 15008 26140
rect 15064 26138 15088 26140
rect 15144 26138 15150 26140
rect 14904 26086 14906 26138
rect 15086 26086 15088 26138
rect 14842 26084 14848 26086
rect 14904 26084 14928 26086
rect 14984 26084 15008 26086
rect 15064 26084 15088 26086
rect 15144 26084 15150 26086
rect 14842 26075 15150 26084
rect 14740 25968 14792 25974
rect 14740 25910 14792 25916
rect 14280 25424 14332 25430
rect 14280 25366 14332 25372
rect 14004 25152 14056 25158
rect 14004 25094 14056 25100
rect 14280 25152 14332 25158
rect 14280 25094 14332 25100
rect 13820 24880 13872 24886
rect 13820 24822 13872 24828
rect 12900 24812 12952 24818
rect 12900 24754 12952 24760
rect 13360 24812 13412 24818
rect 13360 24754 13412 24760
rect 13912 24812 13964 24818
rect 13912 24754 13964 24760
rect 12256 24608 12308 24614
rect 12256 24550 12308 24556
rect 12072 24268 12124 24274
rect 12072 24210 12124 24216
rect 10416 24132 10468 24138
rect 10416 24074 10468 24080
rect 11152 24132 11204 24138
rect 11152 24074 11204 24080
rect 10428 23798 10456 24074
rect 10416 23792 10468 23798
rect 10416 23734 10468 23740
rect 9588 23656 9640 23662
rect 9588 23598 9640 23604
rect 13924 23526 13952 24754
rect 14292 23866 14320 25094
rect 14752 24818 14780 25910
rect 15396 25906 15424 27814
rect 15476 27532 15528 27538
rect 15476 27474 15528 27480
rect 15488 26246 15516 27474
rect 15672 27441 15700 29294
rect 16040 29220 16068 29514
rect 15764 29192 16068 29220
rect 15764 29034 15792 29192
rect 16028 29096 16080 29102
rect 16028 29038 16080 29044
rect 15752 29028 15804 29034
rect 15752 28970 15804 28976
rect 15936 28620 15988 28626
rect 15936 28562 15988 28568
rect 15844 28484 15896 28490
rect 15844 28426 15896 28432
rect 15856 28082 15884 28426
rect 15948 28218 15976 28562
rect 15936 28212 15988 28218
rect 15936 28154 15988 28160
rect 15948 28082 15976 28154
rect 15844 28076 15896 28082
rect 15844 28018 15896 28024
rect 15936 28076 15988 28082
rect 15936 28018 15988 28024
rect 16040 27962 16068 29038
rect 16132 28762 16160 30806
rect 16212 30660 16264 30666
rect 16212 30602 16264 30608
rect 16224 30394 16252 30602
rect 16304 30592 16356 30598
rect 16304 30534 16356 30540
rect 16212 30388 16264 30394
rect 16212 30330 16264 30336
rect 16210 29744 16266 29753
rect 16210 29679 16266 29688
rect 16224 29646 16252 29679
rect 16212 29640 16264 29646
rect 16212 29582 16264 29588
rect 16210 29472 16266 29481
rect 16210 29407 16266 29416
rect 16224 29102 16252 29407
rect 16212 29096 16264 29102
rect 16212 29038 16264 29044
rect 16120 28756 16172 28762
rect 16120 28698 16172 28704
rect 15856 27934 16068 27962
rect 15752 27464 15804 27470
rect 15658 27432 15714 27441
rect 15752 27406 15804 27412
rect 15658 27367 15714 27376
rect 15764 27033 15792 27406
rect 15856 27402 15884 27934
rect 16028 27872 16080 27878
rect 16028 27814 16080 27820
rect 15936 27600 15988 27606
rect 15934 27568 15936 27577
rect 15988 27568 15990 27577
rect 15934 27503 15990 27512
rect 15844 27396 15896 27402
rect 15844 27338 15896 27344
rect 15936 27396 15988 27402
rect 15936 27338 15988 27344
rect 15948 27130 15976 27338
rect 15936 27124 15988 27130
rect 15936 27066 15988 27072
rect 15750 27024 15806 27033
rect 15750 26959 15806 26968
rect 15948 26858 15976 27066
rect 15936 26852 15988 26858
rect 15936 26794 15988 26800
rect 15476 26240 15528 26246
rect 15476 26182 15528 26188
rect 15384 25900 15436 25906
rect 15384 25842 15436 25848
rect 15488 25838 15516 26182
rect 16040 25945 16068 27814
rect 16132 26450 16160 28698
rect 16224 26926 16252 29038
rect 16316 28966 16344 30534
rect 16304 28960 16356 28966
rect 16304 28902 16356 28908
rect 16304 28688 16356 28694
rect 16304 28630 16356 28636
rect 16212 26920 16264 26926
rect 16212 26862 16264 26868
rect 16120 26444 16172 26450
rect 16120 26386 16172 26392
rect 16316 26353 16344 28630
rect 16408 27606 16436 31758
rect 17144 31754 17172 33200
rect 17144 31726 17264 31754
rect 17236 31414 17264 31726
rect 17224 31408 17276 31414
rect 17224 31350 17276 31356
rect 16580 31340 16632 31346
rect 16580 31282 16632 31288
rect 16486 30696 16542 30705
rect 16486 30631 16542 30640
rect 16500 30598 16528 30631
rect 16488 30592 16540 30598
rect 16488 30534 16540 30540
rect 16488 30388 16540 30394
rect 16488 30330 16540 30336
rect 16500 28014 16528 30330
rect 16592 30297 16620 31282
rect 17868 31272 17920 31278
rect 17868 31214 17920 31220
rect 17880 31113 17908 31214
rect 17960 31204 18012 31210
rect 17960 31146 18012 31152
rect 16670 31104 16726 31113
rect 16670 31039 16726 31048
rect 17866 31104 17922 31113
rect 17866 31039 17922 31048
rect 16578 30288 16634 30297
rect 16578 30223 16634 30232
rect 16684 29646 16712 31039
rect 16856 30796 16908 30802
rect 16856 30738 16908 30744
rect 16764 30660 16816 30666
rect 16764 30602 16816 30608
rect 16580 29640 16632 29646
rect 16580 29582 16632 29588
rect 16672 29640 16724 29646
rect 16672 29582 16724 29588
rect 16592 28744 16620 29582
rect 16670 29472 16726 29481
rect 16670 29407 16726 29416
rect 16684 29306 16712 29407
rect 16672 29300 16724 29306
rect 16672 29242 16724 29248
rect 16670 29200 16726 29209
rect 16670 29135 16672 29144
rect 16724 29135 16726 29144
rect 16672 29106 16724 29112
rect 16776 28937 16804 30602
rect 16868 29034 16896 30738
rect 17316 30728 17368 30734
rect 17500 30728 17552 30734
rect 17368 30688 17448 30716
rect 17316 30670 17368 30676
rect 17040 30592 17092 30598
rect 17040 30534 17092 30540
rect 16948 30048 17000 30054
rect 16948 29990 17000 29996
rect 16856 29028 16908 29034
rect 16856 28970 16908 28976
rect 16762 28928 16818 28937
rect 16762 28863 16818 28872
rect 16592 28716 16712 28744
rect 16580 28620 16632 28626
rect 16580 28562 16632 28568
rect 16488 28008 16540 28014
rect 16488 27950 16540 27956
rect 16592 27946 16620 28562
rect 16580 27940 16632 27946
rect 16580 27882 16632 27888
rect 16396 27600 16448 27606
rect 16684 27554 16712 28716
rect 16960 28558 16988 29990
rect 17052 29073 17080 30534
rect 17316 30388 17368 30394
rect 17316 30330 17368 30336
rect 17224 30116 17276 30122
rect 17224 30058 17276 30064
rect 17132 30048 17184 30054
rect 17132 29990 17184 29996
rect 17144 29889 17172 29990
rect 17130 29880 17186 29889
rect 17236 29850 17264 30058
rect 17130 29815 17186 29824
rect 17224 29844 17276 29850
rect 17224 29786 17276 29792
rect 17224 29640 17276 29646
rect 17328 29617 17356 30330
rect 17224 29582 17276 29588
rect 17314 29608 17370 29617
rect 17132 29504 17184 29510
rect 17132 29446 17184 29452
rect 17038 29064 17094 29073
rect 17038 28999 17094 29008
rect 17040 28960 17092 28966
rect 17040 28902 17092 28908
rect 16948 28552 17000 28558
rect 16948 28494 17000 28500
rect 16396 27542 16448 27548
rect 16592 27526 16712 27554
rect 16302 26344 16358 26353
rect 16302 26279 16358 26288
rect 16026 25936 16082 25945
rect 16026 25871 16082 25880
rect 15476 25832 15528 25838
rect 15476 25774 15528 25780
rect 16592 25362 16620 27526
rect 16672 27464 16724 27470
rect 16672 27406 16724 27412
rect 16856 27464 16908 27470
rect 16856 27406 16908 27412
rect 16580 25356 16632 25362
rect 16580 25298 16632 25304
rect 14842 25052 15150 25061
rect 14842 25050 14848 25052
rect 14904 25050 14928 25052
rect 14984 25050 15008 25052
rect 15064 25050 15088 25052
rect 15144 25050 15150 25052
rect 14904 24998 14906 25050
rect 15086 24998 15088 25050
rect 14842 24996 14848 24998
rect 14904 24996 14928 24998
rect 14984 24996 15008 24998
rect 15064 24996 15088 24998
rect 15144 24996 15150 24998
rect 14842 24987 15150 24996
rect 14740 24812 14792 24818
rect 14740 24754 14792 24760
rect 16684 24342 16712 27406
rect 16868 25770 16896 27406
rect 17052 27130 17080 28902
rect 17144 27713 17172 29446
rect 17236 29170 17264 29582
rect 17314 29543 17370 29552
rect 17328 29510 17356 29543
rect 17316 29504 17368 29510
rect 17316 29446 17368 29452
rect 17224 29164 17276 29170
rect 17224 29106 17276 29112
rect 17316 28552 17368 28558
rect 17316 28494 17368 28500
rect 17130 27704 17186 27713
rect 17130 27639 17186 27648
rect 17040 27124 17092 27130
rect 17040 27066 17092 27072
rect 17328 26761 17356 28494
rect 17314 26752 17370 26761
rect 17314 26687 17370 26696
rect 17132 25900 17184 25906
rect 17132 25842 17184 25848
rect 16856 25764 16908 25770
rect 16856 25706 16908 25712
rect 16672 24336 16724 24342
rect 16672 24278 16724 24284
rect 14842 23964 15150 23973
rect 14842 23962 14848 23964
rect 14904 23962 14928 23964
rect 14984 23962 15008 23964
rect 15064 23962 15088 23964
rect 15144 23962 15150 23964
rect 14904 23910 14906 23962
rect 15086 23910 15088 23962
rect 14842 23908 14848 23910
rect 14904 23908 14928 23910
rect 14984 23908 15008 23910
rect 15064 23908 15088 23910
rect 15144 23908 15150 23910
rect 14842 23899 15150 23908
rect 14280 23860 14332 23866
rect 14280 23802 14332 23808
rect 13912 23520 13964 23526
rect 13912 23462 13964 23468
rect 11369 23420 11677 23429
rect 11369 23418 11375 23420
rect 11431 23418 11455 23420
rect 11511 23418 11535 23420
rect 11591 23418 11615 23420
rect 11671 23418 11677 23420
rect 11431 23366 11433 23418
rect 11613 23366 11615 23418
rect 11369 23364 11375 23366
rect 11431 23364 11455 23366
rect 11511 23364 11535 23366
rect 11591 23364 11615 23366
rect 11671 23364 11677 23366
rect 11369 23355 11677 23364
rect 9220 23316 9272 23322
rect 9220 23258 9272 23264
rect 7896 22876 8204 22885
rect 7896 22874 7902 22876
rect 7958 22874 7982 22876
rect 8038 22874 8062 22876
rect 8118 22874 8142 22876
rect 8198 22874 8204 22876
rect 7958 22822 7960 22874
rect 8140 22822 8142 22874
rect 7896 22820 7902 22822
rect 7958 22820 7982 22822
rect 8038 22820 8062 22822
rect 8118 22820 8142 22822
rect 8198 22820 8204 22822
rect 7896 22811 8204 22820
rect 14842 22876 15150 22885
rect 14842 22874 14848 22876
rect 14904 22874 14928 22876
rect 14984 22874 15008 22876
rect 15064 22874 15088 22876
rect 15144 22874 15150 22876
rect 14904 22822 14906 22874
rect 15086 22822 15088 22874
rect 14842 22820 14848 22822
rect 14904 22820 14928 22822
rect 14984 22820 15008 22822
rect 15064 22820 15088 22822
rect 15144 22820 15150 22822
rect 14842 22811 15150 22820
rect 1584 22432 1636 22438
rect 1584 22374 1636 22380
rect 1596 22137 1624 22374
rect 4423 22332 4731 22341
rect 4423 22330 4429 22332
rect 4485 22330 4509 22332
rect 4565 22330 4589 22332
rect 4645 22330 4669 22332
rect 4725 22330 4731 22332
rect 4485 22278 4487 22330
rect 4667 22278 4669 22330
rect 4423 22276 4429 22278
rect 4485 22276 4509 22278
rect 4565 22276 4589 22278
rect 4645 22276 4669 22278
rect 4725 22276 4731 22278
rect 4423 22267 4731 22276
rect 11369 22332 11677 22341
rect 11369 22330 11375 22332
rect 11431 22330 11455 22332
rect 11511 22330 11535 22332
rect 11591 22330 11615 22332
rect 11671 22330 11677 22332
rect 11431 22278 11433 22330
rect 11613 22278 11615 22330
rect 11369 22276 11375 22278
rect 11431 22276 11455 22278
rect 11511 22276 11535 22278
rect 11591 22276 11615 22278
rect 11671 22276 11677 22278
rect 11369 22267 11677 22276
rect 1582 22128 1638 22137
rect 1582 22063 1638 22072
rect 7896 21788 8204 21797
rect 7896 21786 7902 21788
rect 7958 21786 7982 21788
rect 8038 21786 8062 21788
rect 8118 21786 8142 21788
rect 8198 21786 8204 21788
rect 7958 21734 7960 21786
rect 8140 21734 8142 21786
rect 7896 21732 7902 21734
rect 7958 21732 7982 21734
rect 8038 21732 8062 21734
rect 8118 21732 8142 21734
rect 8198 21732 8204 21734
rect 7896 21723 8204 21732
rect 14842 21788 15150 21797
rect 14842 21786 14848 21788
rect 14904 21786 14928 21788
rect 14984 21786 15008 21788
rect 15064 21786 15088 21788
rect 15144 21786 15150 21788
rect 14904 21734 14906 21786
rect 15086 21734 15088 21786
rect 14842 21732 14848 21734
rect 14904 21732 14928 21734
rect 14984 21732 15008 21734
rect 15064 21732 15088 21734
rect 15144 21732 15150 21734
rect 14842 21723 15150 21732
rect 1584 21480 1636 21486
rect 1582 21448 1584 21457
rect 1636 21448 1638 21457
rect 1582 21383 1638 21392
rect 4423 21244 4731 21253
rect 4423 21242 4429 21244
rect 4485 21242 4509 21244
rect 4565 21242 4589 21244
rect 4645 21242 4669 21244
rect 4725 21242 4731 21244
rect 4485 21190 4487 21242
rect 4667 21190 4669 21242
rect 4423 21188 4429 21190
rect 4485 21188 4509 21190
rect 4565 21188 4589 21190
rect 4645 21188 4669 21190
rect 4725 21188 4731 21190
rect 4423 21179 4731 21188
rect 11369 21244 11677 21253
rect 11369 21242 11375 21244
rect 11431 21242 11455 21244
rect 11511 21242 11535 21244
rect 11591 21242 11615 21244
rect 11671 21242 11677 21244
rect 11431 21190 11433 21242
rect 11613 21190 11615 21242
rect 11369 21188 11375 21190
rect 11431 21188 11455 21190
rect 11511 21188 11535 21190
rect 11591 21188 11615 21190
rect 11671 21188 11677 21190
rect 11369 21179 11677 21188
rect 7896 20700 8204 20709
rect 7896 20698 7902 20700
rect 7958 20698 7982 20700
rect 8038 20698 8062 20700
rect 8118 20698 8142 20700
rect 8198 20698 8204 20700
rect 7958 20646 7960 20698
rect 8140 20646 8142 20698
rect 7896 20644 7902 20646
rect 7958 20644 7982 20646
rect 8038 20644 8062 20646
rect 8118 20644 8142 20646
rect 8198 20644 8204 20646
rect 7896 20635 8204 20644
rect 14842 20700 15150 20709
rect 14842 20698 14848 20700
rect 14904 20698 14928 20700
rect 14984 20698 15008 20700
rect 15064 20698 15088 20700
rect 15144 20698 15150 20700
rect 14904 20646 14906 20698
rect 15086 20646 15088 20698
rect 14842 20644 14848 20646
rect 14904 20644 14928 20646
rect 14984 20644 15008 20646
rect 15064 20644 15088 20646
rect 15144 20644 15150 20646
rect 14842 20635 15150 20644
rect 1584 20256 1636 20262
rect 1584 20198 1636 20204
rect 1596 20097 1624 20198
rect 4423 20156 4731 20165
rect 4423 20154 4429 20156
rect 4485 20154 4509 20156
rect 4565 20154 4589 20156
rect 4645 20154 4669 20156
rect 4725 20154 4731 20156
rect 4485 20102 4487 20154
rect 4667 20102 4669 20154
rect 4423 20100 4429 20102
rect 4485 20100 4509 20102
rect 4565 20100 4589 20102
rect 4645 20100 4669 20102
rect 4725 20100 4731 20102
rect 1582 20088 1638 20097
rect 4423 20091 4731 20100
rect 11369 20156 11677 20165
rect 11369 20154 11375 20156
rect 11431 20154 11455 20156
rect 11511 20154 11535 20156
rect 11591 20154 11615 20156
rect 11671 20154 11677 20156
rect 11431 20102 11433 20154
rect 11613 20102 11615 20154
rect 11369 20100 11375 20102
rect 11431 20100 11455 20102
rect 11511 20100 11535 20102
rect 11591 20100 11615 20102
rect 11671 20100 11677 20102
rect 11369 20091 11677 20100
rect 1582 20023 1638 20032
rect 1584 19848 1636 19854
rect 1584 19790 1636 19796
rect 1596 19417 1624 19790
rect 7896 19612 8204 19621
rect 7896 19610 7902 19612
rect 7958 19610 7982 19612
rect 8038 19610 8062 19612
rect 8118 19610 8142 19612
rect 8198 19610 8204 19612
rect 7958 19558 7960 19610
rect 8140 19558 8142 19610
rect 7896 19556 7902 19558
rect 7958 19556 7982 19558
rect 8038 19556 8062 19558
rect 8118 19556 8142 19558
rect 8198 19556 8204 19558
rect 7896 19547 8204 19556
rect 14842 19612 15150 19621
rect 14842 19610 14848 19612
rect 14904 19610 14928 19612
rect 14984 19610 15008 19612
rect 15064 19610 15088 19612
rect 15144 19610 15150 19612
rect 14904 19558 14906 19610
rect 15086 19558 15088 19610
rect 14842 19556 14848 19558
rect 14904 19556 14928 19558
rect 14984 19556 15008 19558
rect 15064 19556 15088 19558
rect 15144 19556 15150 19558
rect 14842 19547 15150 19556
rect 1582 19408 1638 19417
rect 1582 19343 1638 19352
rect 4423 19068 4731 19077
rect 4423 19066 4429 19068
rect 4485 19066 4509 19068
rect 4565 19066 4589 19068
rect 4645 19066 4669 19068
rect 4725 19066 4731 19068
rect 4485 19014 4487 19066
rect 4667 19014 4669 19066
rect 4423 19012 4429 19014
rect 4485 19012 4509 19014
rect 4565 19012 4589 19014
rect 4645 19012 4669 19014
rect 4725 19012 4731 19014
rect 4423 19003 4731 19012
rect 11369 19068 11677 19077
rect 11369 19066 11375 19068
rect 11431 19066 11455 19068
rect 11511 19066 11535 19068
rect 11591 19066 11615 19068
rect 11671 19066 11677 19068
rect 11431 19014 11433 19066
rect 11613 19014 11615 19066
rect 11369 19012 11375 19014
rect 11431 19012 11455 19014
rect 11511 19012 11535 19014
rect 11591 19012 11615 19014
rect 11671 19012 11677 19014
rect 11369 19003 11677 19012
rect 7896 18524 8204 18533
rect 7896 18522 7902 18524
rect 7958 18522 7982 18524
rect 8038 18522 8062 18524
rect 8118 18522 8142 18524
rect 8198 18522 8204 18524
rect 7958 18470 7960 18522
rect 8140 18470 8142 18522
rect 7896 18468 7902 18470
rect 7958 18468 7982 18470
rect 8038 18468 8062 18470
rect 8118 18468 8142 18470
rect 8198 18468 8204 18470
rect 7896 18459 8204 18468
rect 14842 18524 15150 18533
rect 14842 18522 14848 18524
rect 14904 18522 14928 18524
rect 14984 18522 15008 18524
rect 15064 18522 15088 18524
rect 15144 18522 15150 18524
rect 14904 18470 14906 18522
rect 15086 18470 15088 18522
rect 14842 18468 14848 18470
rect 14904 18468 14928 18470
rect 14984 18468 15008 18470
rect 15064 18468 15088 18470
rect 15144 18468 15150 18470
rect 14842 18459 15150 18468
rect 1584 18080 1636 18086
rect 1582 18048 1584 18057
rect 1636 18048 1638 18057
rect 1582 17983 1638 17992
rect 4423 17980 4731 17989
rect 4423 17978 4429 17980
rect 4485 17978 4509 17980
rect 4565 17978 4589 17980
rect 4645 17978 4669 17980
rect 4725 17978 4731 17980
rect 4485 17926 4487 17978
rect 4667 17926 4669 17978
rect 4423 17924 4429 17926
rect 4485 17924 4509 17926
rect 4565 17924 4589 17926
rect 4645 17924 4669 17926
rect 4725 17924 4731 17926
rect 4423 17915 4731 17924
rect 11369 17980 11677 17989
rect 11369 17978 11375 17980
rect 11431 17978 11455 17980
rect 11511 17978 11535 17980
rect 11591 17978 11615 17980
rect 11671 17978 11677 17980
rect 11431 17926 11433 17978
rect 11613 17926 11615 17978
rect 11369 17924 11375 17926
rect 11431 17924 11455 17926
rect 11511 17924 11535 17926
rect 11591 17924 11615 17926
rect 11671 17924 11677 17926
rect 11369 17915 11677 17924
rect 1584 17672 1636 17678
rect 1584 17614 1636 17620
rect 1596 17377 1624 17614
rect 7896 17436 8204 17445
rect 7896 17434 7902 17436
rect 7958 17434 7982 17436
rect 8038 17434 8062 17436
rect 8118 17434 8142 17436
rect 8198 17434 8204 17436
rect 7958 17382 7960 17434
rect 8140 17382 8142 17434
rect 7896 17380 7902 17382
rect 7958 17380 7982 17382
rect 8038 17380 8062 17382
rect 8118 17380 8142 17382
rect 8198 17380 8204 17382
rect 1582 17368 1638 17377
rect 7896 17371 8204 17380
rect 14842 17436 15150 17445
rect 14842 17434 14848 17436
rect 14904 17434 14928 17436
rect 14984 17434 15008 17436
rect 15064 17434 15088 17436
rect 15144 17434 15150 17436
rect 14904 17382 14906 17434
rect 15086 17382 15088 17434
rect 14842 17380 14848 17382
rect 14904 17380 14928 17382
rect 14984 17380 15008 17382
rect 15064 17380 15088 17382
rect 15144 17380 15150 17382
rect 14842 17371 15150 17380
rect 1582 17303 1638 17312
rect 4423 16892 4731 16901
rect 4423 16890 4429 16892
rect 4485 16890 4509 16892
rect 4565 16890 4589 16892
rect 4645 16890 4669 16892
rect 4725 16890 4731 16892
rect 4485 16838 4487 16890
rect 4667 16838 4669 16890
rect 4423 16836 4429 16838
rect 4485 16836 4509 16838
rect 4565 16836 4589 16838
rect 4645 16836 4669 16838
rect 4725 16836 4731 16838
rect 4423 16827 4731 16836
rect 11369 16892 11677 16901
rect 11369 16890 11375 16892
rect 11431 16890 11455 16892
rect 11511 16890 11535 16892
rect 11591 16890 11615 16892
rect 11671 16890 11677 16892
rect 11431 16838 11433 16890
rect 11613 16838 11615 16890
rect 11369 16836 11375 16838
rect 11431 16836 11455 16838
rect 11511 16836 11535 16838
rect 11591 16836 11615 16838
rect 11671 16836 11677 16838
rect 11369 16827 11677 16836
rect 7896 16348 8204 16357
rect 7896 16346 7902 16348
rect 7958 16346 7982 16348
rect 8038 16346 8062 16348
rect 8118 16346 8142 16348
rect 8198 16346 8204 16348
rect 7958 16294 7960 16346
rect 8140 16294 8142 16346
rect 7896 16292 7902 16294
rect 7958 16292 7982 16294
rect 8038 16292 8062 16294
rect 8118 16292 8142 16294
rect 8198 16292 8204 16294
rect 7896 16283 8204 16292
rect 14842 16348 15150 16357
rect 14842 16346 14848 16348
rect 14904 16346 14928 16348
rect 14984 16346 15008 16348
rect 15064 16346 15088 16348
rect 15144 16346 15150 16348
rect 14904 16294 14906 16346
rect 15086 16294 15088 16346
rect 14842 16292 14848 16294
rect 14904 16292 14928 16294
rect 14984 16292 15008 16294
rect 15064 16292 15088 16294
rect 15144 16292 15150 16294
rect 14842 16283 15150 16292
rect 1584 16040 1636 16046
rect 1582 16008 1584 16017
rect 1636 16008 1638 16017
rect 1582 15943 1638 15952
rect 4423 15804 4731 15813
rect 4423 15802 4429 15804
rect 4485 15802 4509 15804
rect 4565 15802 4589 15804
rect 4645 15802 4669 15804
rect 4725 15802 4731 15804
rect 4485 15750 4487 15802
rect 4667 15750 4669 15802
rect 4423 15748 4429 15750
rect 4485 15748 4509 15750
rect 4565 15748 4589 15750
rect 4645 15748 4669 15750
rect 4725 15748 4731 15750
rect 4423 15739 4731 15748
rect 11369 15804 11677 15813
rect 11369 15802 11375 15804
rect 11431 15802 11455 15804
rect 11511 15802 11535 15804
rect 11591 15802 11615 15804
rect 11671 15802 11677 15804
rect 11431 15750 11433 15802
rect 11613 15750 11615 15802
rect 11369 15748 11375 15750
rect 11431 15748 11455 15750
rect 11511 15748 11535 15750
rect 11591 15748 11615 15750
rect 11671 15748 11677 15750
rect 11369 15739 11677 15748
rect 1584 15496 1636 15502
rect 1584 15438 1636 15444
rect 1596 15337 1624 15438
rect 1582 15328 1638 15337
rect 1582 15263 1638 15272
rect 7896 15260 8204 15269
rect 7896 15258 7902 15260
rect 7958 15258 7982 15260
rect 8038 15258 8062 15260
rect 8118 15258 8142 15260
rect 8198 15258 8204 15260
rect 7958 15206 7960 15258
rect 8140 15206 8142 15258
rect 7896 15204 7902 15206
rect 7958 15204 7982 15206
rect 8038 15204 8062 15206
rect 8118 15204 8142 15206
rect 8198 15204 8204 15206
rect 7896 15195 8204 15204
rect 14842 15260 15150 15269
rect 14842 15258 14848 15260
rect 14904 15258 14928 15260
rect 14984 15258 15008 15260
rect 15064 15258 15088 15260
rect 15144 15258 15150 15260
rect 14904 15206 14906 15258
rect 15086 15206 15088 15258
rect 14842 15204 14848 15206
rect 14904 15204 14928 15206
rect 14984 15204 15008 15206
rect 15064 15204 15088 15206
rect 15144 15204 15150 15206
rect 14842 15195 15150 15204
rect 4423 14716 4731 14725
rect 4423 14714 4429 14716
rect 4485 14714 4509 14716
rect 4565 14714 4589 14716
rect 4645 14714 4669 14716
rect 4725 14714 4731 14716
rect 4485 14662 4487 14714
rect 4667 14662 4669 14714
rect 4423 14660 4429 14662
rect 4485 14660 4509 14662
rect 4565 14660 4589 14662
rect 4645 14660 4669 14662
rect 4725 14660 4731 14662
rect 4423 14651 4731 14660
rect 11369 14716 11677 14725
rect 11369 14714 11375 14716
rect 11431 14714 11455 14716
rect 11511 14714 11535 14716
rect 11591 14714 11615 14716
rect 11671 14714 11677 14716
rect 11431 14662 11433 14714
rect 11613 14662 11615 14714
rect 11369 14660 11375 14662
rect 11431 14660 11455 14662
rect 11511 14660 11535 14662
rect 11591 14660 11615 14662
rect 11671 14660 11677 14662
rect 11369 14651 11677 14660
rect 1584 14408 1636 14414
rect 1584 14350 1636 14356
rect 1596 13977 1624 14350
rect 7896 14172 8204 14181
rect 7896 14170 7902 14172
rect 7958 14170 7982 14172
rect 8038 14170 8062 14172
rect 8118 14170 8142 14172
rect 8198 14170 8204 14172
rect 7958 14118 7960 14170
rect 8140 14118 8142 14170
rect 7896 14116 7902 14118
rect 7958 14116 7982 14118
rect 8038 14116 8062 14118
rect 8118 14116 8142 14118
rect 8198 14116 8204 14118
rect 7896 14107 8204 14116
rect 14842 14172 15150 14181
rect 14842 14170 14848 14172
rect 14904 14170 14928 14172
rect 14984 14170 15008 14172
rect 15064 14170 15088 14172
rect 15144 14170 15150 14172
rect 14904 14118 14906 14170
rect 15086 14118 15088 14170
rect 14842 14116 14848 14118
rect 14904 14116 14928 14118
rect 14984 14116 15008 14118
rect 15064 14116 15088 14118
rect 15144 14116 15150 14118
rect 14842 14107 15150 14116
rect 1582 13968 1638 13977
rect 1582 13903 1638 13912
rect 4423 13628 4731 13637
rect 4423 13626 4429 13628
rect 4485 13626 4509 13628
rect 4565 13626 4589 13628
rect 4645 13626 4669 13628
rect 4725 13626 4731 13628
rect 4485 13574 4487 13626
rect 4667 13574 4669 13626
rect 4423 13572 4429 13574
rect 4485 13572 4509 13574
rect 4565 13572 4589 13574
rect 4645 13572 4669 13574
rect 4725 13572 4731 13574
rect 4423 13563 4731 13572
rect 11369 13628 11677 13637
rect 11369 13626 11375 13628
rect 11431 13626 11455 13628
rect 11511 13626 11535 13628
rect 11591 13626 11615 13628
rect 11671 13626 11677 13628
rect 11431 13574 11433 13626
rect 11613 13574 11615 13626
rect 11369 13572 11375 13574
rect 11431 13572 11455 13574
rect 11511 13572 11535 13574
rect 11591 13572 11615 13574
rect 11671 13572 11677 13574
rect 11369 13563 11677 13572
rect 1584 13320 1636 13326
rect 1582 13288 1584 13297
rect 1636 13288 1638 13297
rect 1582 13223 1638 13232
rect 7896 13084 8204 13093
rect 7896 13082 7902 13084
rect 7958 13082 7982 13084
rect 8038 13082 8062 13084
rect 8118 13082 8142 13084
rect 8198 13082 8204 13084
rect 7958 13030 7960 13082
rect 8140 13030 8142 13082
rect 7896 13028 7902 13030
rect 7958 13028 7982 13030
rect 8038 13028 8062 13030
rect 8118 13028 8142 13030
rect 8198 13028 8204 13030
rect 7896 13019 8204 13028
rect 14842 13084 15150 13093
rect 14842 13082 14848 13084
rect 14904 13082 14928 13084
rect 14984 13082 15008 13084
rect 15064 13082 15088 13084
rect 15144 13082 15150 13084
rect 14904 13030 14906 13082
rect 15086 13030 15088 13082
rect 14842 13028 14848 13030
rect 14904 13028 14928 13030
rect 14984 13028 15008 13030
rect 15064 13028 15088 13030
rect 15144 13028 15150 13030
rect 14842 13019 15150 13028
rect 4423 12540 4731 12549
rect 4423 12538 4429 12540
rect 4485 12538 4509 12540
rect 4565 12538 4589 12540
rect 4645 12538 4669 12540
rect 4725 12538 4731 12540
rect 4485 12486 4487 12538
rect 4667 12486 4669 12538
rect 4423 12484 4429 12486
rect 4485 12484 4509 12486
rect 4565 12484 4589 12486
rect 4645 12484 4669 12486
rect 4725 12484 4731 12486
rect 4423 12475 4731 12484
rect 11369 12540 11677 12549
rect 11369 12538 11375 12540
rect 11431 12538 11455 12540
rect 11511 12538 11535 12540
rect 11591 12538 11615 12540
rect 11671 12538 11677 12540
rect 11431 12486 11433 12538
rect 11613 12486 11615 12538
rect 11369 12484 11375 12486
rect 11431 12484 11455 12486
rect 11511 12484 11535 12486
rect 11591 12484 11615 12486
rect 11671 12484 11677 12486
rect 11369 12475 11677 12484
rect 1584 12232 1636 12238
rect 1584 12174 1636 12180
rect 1596 11937 1624 12174
rect 7896 11996 8204 12005
rect 7896 11994 7902 11996
rect 7958 11994 7982 11996
rect 8038 11994 8062 11996
rect 8118 11994 8142 11996
rect 8198 11994 8204 11996
rect 7958 11942 7960 11994
rect 8140 11942 8142 11994
rect 7896 11940 7902 11942
rect 7958 11940 7982 11942
rect 8038 11940 8062 11942
rect 8118 11940 8142 11942
rect 8198 11940 8204 11942
rect 1582 11928 1638 11937
rect 7896 11931 8204 11940
rect 14842 11996 15150 12005
rect 14842 11994 14848 11996
rect 14904 11994 14928 11996
rect 14984 11994 15008 11996
rect 15064 11994 15088 11996
rect 15144 11994 15150 11996
rect 14904 11942 14906 11994
rect 15086 11942 15088 11994
rect 14842 11940 14848 11942
rect 14904 11940 14928 11942
rect 14984 11940 15008 11942
rect 15064 11940 15088 11942
rect 15144 11940 15150 11942
rect 14842 11931 15150 11940
rect 1582 11863 1638 11872
rect 1584 11552 1636 11558
rect 1584 11494 1636 11500
rect 1596 11257 1624 11494
rect 4423 11452 4731 11461
rect 4423 11450 4429 11452
rect 4485 11450 4509 11452
rect 4565 11450 4589 11452
rect 4645 11450 4669 11452
rect 4725 11450 4731 11452
rect 4485 11398 4487 11450
rect 4667 11398 4669 11450
rect 4423 11396 4429 11398
rect 4485 11396 4509 11398
rect 4565 11396 4589 11398
rect 4645 11396 4669 11398
rect 4725 11396 4731 11398
rect 4423 11387 4731 11396
rect 11369 11452 11677 11461
rect 11369 11450 11375 11452
rect 11431 11450 11455 11452
rect 11511 11450 11535 11452
rect 11591 11450 11615 11452
rect 11671 11450 11677 11452
rect 11431 11398 11433 11450
rect 11613 11398 11615 11450
rect 11369 11396 11375 11398
rect 11431 11396 11455 11398
rect 11511 11396 11535 11398
rect 11591 11396 11615 11398
rect 11671 11396 11677 11398
rect 11369 11387 11677 11396
rect 1582 11248 1638 11257
rect 1582 11183 1638 11192
rect 7896 10908 8204 10917
rect 7896 10906 7902 10908
rect 7958 10906 7982 10908
rect 8038 10906 8062 10908
rect 8118 10906 8142 10908
rect 8198 10906 8204 10908
rect 7958 10854 7960 10906
rect 8140 10854 8142 10906
rect 7896 10852 7902 10854
rect 7958 10852 7982 10854
rect 8038 10852 8062 10854
rect 8118 10852 8142 10854
rect 8198 10852 8204 10854
rect 7896 10843 8204 10852
rect 14842 10908 15150 10917
rect 14842 10906 14848 10908
rect 14904 10906 14928 10908
rect 14984 10906 15008 10908
rect 15064 10906 15088 10908
rect 15144 10906 15150 10908
rect 14904 10854 14906 10906
rect 15086 10854 15088 10906
rect 14842 10852 14848 10854
rect 14904 10852 14928 10854
rect 14984 10852 15008 10854
rect 15064 10852 15088 10854
rect 15144 10852 15150 10854
rect 14842 10843 15150 10852
rect 4423 10364 4731 10373
rect 4423 10362 4429 10364
rect 4485 10362 4509 10364
rect 4565 10362 4589 10364
rect 4645 10362 4669 10364
rect 4725 10362 4731 10364
rect 4485 10310 4487 10362
rect 4667 10310 4669 10362
rect 4423 10308 4429 10310
rect 4485 10308 4509 10310
rect 4565 10308 4589 10310
rect 4645 10308 4669 10310
rect 4725 10308 4731 10310
rect 4423 10299 4731 10308
rect 11369 10364 11677 10373
rect 11369 10362 11375 10364
rect 11431 10362 11455 10364
rect 11511 10362 11535 10364
rect 11591 10362 11615 10364
rect 11671 10362 11677 10364
rect 11431 10310 11433 10362
rect 11613 10310 11615 10362
rect 11369 10308 11375 10310
rect 11431 10308 11455 10310
rect 11511 10308 11535 10310
rect 11591 10308 11615 10310
rect 11671 10308 11677 10310
rect 11369 10299 11677 10308
rect 1584 10056 1636 10062
rect 1584 9998 1636 10004
rect 1596 9897 1624 9998
rect 1582 9888 1638 9897
rect 1582 9823 1638 9832
rect 7896 9820 8204 9829
rect 7896 9818 7902 9820
rect 7958 9818 7982 9820
rect 8038 9818 8062 9820
rect 8118 9818 8142 9820
rect 8198 9818 8204 9820
rect 7958 9766 7960 9818
rect 8140 9766 8142 9818
rect 7896 9764 7902 9766
rect 7958 9764 7982 9766
rect 8038 9764 8062 9766
rect 8118 9764 8142 9766
rect 8198 9764 8204 9766
rect 7896 9755 8204 9764
rect 14842 9820 15150 9829
rect 14842 9818 14848 9820
rect 14904 9818 14928 9820
rect 14984 9818 15008 9820
rect 15064 9818 15088 9820
rect 15144 9818 15150 9820
rect 14904 9766 14906 9818
rect 15086 9766 15088 9818
rect 14842 9764 14848 9766
rect 14904 9764 14928 9766
rect 14984 9764 15008 9766
rect 15064 9764 15088 9766
rect 15144 9764 15150 9766
rect 14842 9755 15150 9764
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1596 9217 1624 9318
rect 4423 9276 4731 9285
rect 4423 9274 4429 9276
rect 4485 9274 4509 9276
rect 4565 9274 4589 9276
rect 4645 9274 4669 9276
rect 4725 9274 4731 9276
rect 4485 9222 4487 9274
rect 4667 9222 4669 9274
rect 4423 9220 4429 9222
rect 4485 9220 4509 9222
rect 4565 9220 4589 9222
rect 4645 9220 4669 9222
rect 4725 9220 4731 9222
rect 1582 9208 1638 9217
rect 4423 9211 4731 9220
rect 11369 9276 11677 9285
rect 11369 9274 11375 9276
rect 11431 9274 11455 9276
rect 11511 9274 11535 9276
rect 11591 9274 11615 9276
rect 11671 9274 11677 9276
rect 11431 9222 11433 9274
rect 11613 9222 11615 9274
rect 11369 9220 11375 9222
rect 11431 9220 11455 9222
rect 11511 9220 11535 9222
rect 11591 9220 11615 9222
rect 11671 9220 11677 9222
rect 11369 9211 11677 9220
rect 1582 9143 1638 9152
rect 7896 8732 8204 8741
rect 7896 8730 7902 8732
rect 7958 8730 7982 8732
rect 8038 8730 8062 8732
rect 8118 8730 8142 8732
rect 8198 8730 8204 8732
rect 7958 8678 7960 8730
rect 8140 8678 8142 8730
rect 7896 8676 7902 8678
rect 7958 8676 7982 8678
rect 8038 8676 8062 8678
rect 8118 8676 8142 8678
rect 8198 8676 8204 8678
rect 7896 8667 8204 8676
rect 14842 8732 15150 8741
rect 14842 8730 14848 8732
rect 14904 8730 14928 8732
rect 14984 8730 15008 8732
rect 15064 8730 15088 8732
rect 15144 8730 15150 8732
rect 14904 8678 14906 8730
rect 15086 8678 15088 8730
rect 14842 8676 14848 8678
rect 14904 8676 14928 8678
rect 14984 8676 15008 8678
rect 15064 8676 15088 8678
rect 15144 8676 15150 8678
rect 14842 8667 15150 8676
rect 4423 8188 4731 8197
rect 4423 8186 4429 8188
rect 4485 8186 4509 8188
rect 4565 8186 4589 8188
rect 4645 8186 4669 8188
rect 4725 8186 4731 8188
rect 4485 8134 4487 8186
rect 4667 8134 4669 8186
rect 4423 8132 4429 8134
rect 4485 8132 4509 8134
rect 4565 8132 4589 8134
rect 4645 8132 4669 8134
rect 4725 8132 4731 8134
rect 4423 8123 4731 8132
rect 11369 8188 11677 8197
rect 11369 8186 11375 8188
rect 11431 8186 11455 8188
rect 11511 8186 11535 8188
rect 11591 8186 11615 8188
rect 11671 8186 11677 8188
rect 11431 8134 11433 8186
rect 11613 8134 11615 8186
rect 11369 8132 11375 8134
rect 11431 8132 11455 8134
rect 11511 8132 11535 8134
rect 11591 8132 11615 8134
rect 11671 8132 11677 8134
rect 11369 8123 11677 8132
rect 1584 7880 1636 7886
rect 1582 7848 1584 7857
rect 1636 7848 1638 7857
rect 1582 7783 1638 7792
rect 7896 7644 8204 7653
rect 7896 7642 7902 7644
rect 7958 7642 7982 7644
rect 8038 7642 8062 7644
rect 8118 7642 8142 7644
rect 8198 7642 8204 7644
rect 7958 7590 7960 7642
rect 8140 7590 8142 7642
rect 7896 7588 7902 7590
rect 7958 7588 7982 7590
rect 8038 7588 8062 7590
rect 8118 7588 8142 7590
rect 8198 7588 8204 7590
rect 7896 7579 8204 7588
rect 14842 7644 15150 7653
rect 14842 7642 14848 7644
rect 14904 7642 14928 7644
rect 14984 7642 15008 7644
rect 15064 7642 15088 7644
rect 15144 7642 15150 7644
rect 14904 7590 14906 7642
rect 15086 7590 15088 7642
rect 14842 7588 14848 7590
rect 14904 7588 14928 7590
rect 14984 7588 15008 7590
rect 15064 7588 15088 7590
rect 15144 7588 15150 7590
rect 14842 7579 15150 7588
rect 1584 7200 1636 7206
rect 1582 7168 1584 7177
rect 1636 7168 1638 7177
rect 1582 7103 1638 7112
rect 4423 7100 4731 7109
rect 4423 7098 4429 7100
rect 4485 7098 4509 7100
rect 4565 7098 4589 7100
rect 4645 7098 4669 7100
rect 4725 7098 4731 7100
rect 4485 7046 4487 7098
rect 4667 7046 4669 7098
rect 4423 7044 4429 7046
rect 4485 7044 4509 7046
rect 4565 7044 4589 7046
rect 4645 7044 4669 7046
rect 4725 7044 4731 7046
rect 4423 7035 4731 7044
rect 11369 7100 11677 7109
rect 11369 7098 11375 7100
rect 11431 7098 11455 7100
rect 11511 7098 11535 7100
rect 11591 7098 11615 7100
rect 11671 7098 11677 7100
rect 11431 7046 11433 7098
rect 11613 7046 11615 7098
rect 11369 7044 11375 7046
rect 11431 7044 11455 7046
rect 11511 7044 11535 7046
rect 11591 7044 11615 7046
rect 11671 7044 11677 7046
rect 11369 7035 11677 7044
rect 7896 6556 8204 6565
rect 7896 6554 7902 6556
rect 7958 6554 7982 6556
rect 8038 6554 8062 6556
rect 8118 6554 8142 6556
rect 8198 6554 8204 6556
rect 7958 6502 7960 6554
rect 8140 6502 8142 6554
rect 7896 6500 7902 6502
rect 7958 6500 7982 6502
rect 8038 6500 8062 6502
rect 8118 6500 8142 6502
rect 8198 6500 8204 6502
rect 7896 6491 8204 6500
rect 14842 6556 15150 6565
rect 14842 6554 14848 6556
rect 14904 6554 14928 6556
rect 14984 6554 15008 6556
rect 15064 6554 15088 6556
rect 15144 6554 15150 6556
rect 14904 6502 14906 6554
rect 15086 6502 15088 6554
rect 14842 6500 14848 6502
rect 14904 6500 14928 6502
rect 14984 6500 15008 6502
rect 15064 6500 15088 6502
rect 15144 6500 15150 6502
rect 14842 6491 15150 6500
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1596 5817 1624 6054
rect 4423 6012 4731 6021
rect 4423 6010 4429 6012
rect 4485 6010 4509 6012
rect 4565 6010 4589 6012
rect 4645 6010 4669 6012
rect 4725 6010 4731 6012
rect 4485 5958 4487 6010
rect 4667 5958 4669 6010
rect 4423 5956 4429 5958
rect 4485 5956 4509 5958
rect 4565 5956 4589 5958
rect 4645 5956 4669 5958
rect 4725 5956 4731 5958
rect 4423 5947 4731 5956
rect 11369 6012 11677 6021
rect 11369 6010 11375 6012
rect 11431 6010 11455 6012
rect 11511 6010 11535 6012
rect 11591 6010 11615 6012
rect 11671 6010 11677 6012
rect 11431 5958 11433 6010
rect 11613 5958 11615 6010
rect 11369 5956 11375 5958
rect 11431 5956 11455 5958
rect 11511 5956 11535 5958
rect 11591 5956 11615 5958
rect 11671 5956 11677 5958
rect 11369 5947 11677 5956
rect 1582 5808 1638 5817
rect 1582 5743 1638 5752
rect 7896 5468 8204 5477
rect 7896 5466 7902 5468
rect 7958 5466 7982 5468
rect 8038 5466 8062 5468
rect 8118 5466 8142 5468
rect 8198 5466 8204 5468
rect 7958 5414 7960 5466
rect 8140 5414 8142 5466
rect 7896 5412 7902 5414
rect 7958 5412 7982 5414
rect 8038 5412 8062 5414
rect 8118 5412 8142 5414
rect 8198 5412 8204 5414
rect 7896 5403 8204 5412
rect 14842 5468 15150 5477
rect 14842 5466 14848 5468
rect 14904 5466 14928 5468
rect 14984 5466 15008 5468
rect 15064 5466 15088 5468
rect 15144 5466 15150 5468
rect 14904 5414 14906 5466
rect 15086 5414 15088 5466
rect 14842 5412 14848 5414
rect 14904 5412 14928 5414
rect 14984 5412 15008 5414
rect 15064 5412 15088 5414
rect 15144 5412 15150 5414
rect 14842 5403 15150 5412
rect 1584 5160 1636 5166
rect 1582 5128 1584 5137
rect 1636 5128 1638 5137
rect 1582 5063 1638 5072
rect 4423 4924 4731 4933
rect 4423 4922 4429 4924
rect 4485 4922 4509 4924
rect 4565 4922 4589 4924
rect 4645 4922 4669 4924
rect 4725 4922 4731 4924
rect 4485 4870 4487 4922
rect 4667 4870 4669 4922
rect 4423 4868 4429 4870
rect 4485 4868 4509 4870
rect 4565 4868 4589 4870
rect 4645 4868 4669 4870
rect 4725 4868 4731 4870
rect 4423 4859 4731 4868
rect 11369 4924 11677 4933
rect 11369 4922 11375 4924
rect 11431 4922 11455 4924
rect 11511 4922 11535 4924
rect 11591 4922 11615 4924
rect 11671 4922 11677 4924
rect 11431 4870 11433 4922
rect 11613 4870 11615 4922
rect 11369 4868 11375 4870
rect 11431 4868 11455 4870
rect 11511 4868 11535 4870
rect 11591 4868 11615 4870
rect 11671 4868 11677 4870
rect 11369 4859 11677 4868
rect 7896 4380 8204 4389
rect 7896 4378 7902 4380
rect 7958 4378 7982 4380
rect 8038 4378 8062 4380
rect 8118 4378 8142 4380
rect 8198 4378 8204 4380
rect 7958 4326 7960 4378
rect 8140 4326 8142 4378
rect 7896 4324 7902 4326
rect 7958 4324 7982 4326
rect 8038 4324 8062 4326
rect 8118 4324 8142 4326
rect 8198 4324 8204 4326
rect 7896 4315 8204 4324
rect 14842 4380 15150 4389
rect 14842 4378 14848 4380
rect 14904 4378 14928 4380
rect 14984 4378 15008 4380
rect 15064 4378 15088 4380
rect 15144 4378 15150 4380
rect 14904 4326 14906 4378
rect 15086 4326 15088 4378
rect 14842 4324 14848 4326
rect 14904 4324 14928 4326
rect 14984 4324 15008 4326
rect 15064 4324 15088 4326
rect 15144 4324 15150 4326
rect 14842 4315 15150 4324
rect 17144 4078 17172 25842
rect 17420 25702 17448 30688
rect 17500 30670 17552 30676
rect 17512 30394 17540 30670
rect 17500 30388 17552 30394
rect 17500 30330 17552 30336
rect 17684 30388 17736 30394
rect 17684 30330 17736 30336
rect 17592 30184 17644 30190
rect 17592 30126 17644 30132
rect 17500 30048 17552 30054
rect 17500 29990 17552 29996
rect 17512 29170 17540 29990
rect 17604 29578 17632 30126
rect 17592 29572 17644 29578
rect 17592 29514 17644 29520
rect 17500 29164 17552 29170
rect 17500 29106 17552 29112
rect 17512 26625 17540 29106
rect 17592 29028 17644 29034
rect 17592 28970 17644 28976
rect 17498 26616 17554 26625
rect 17498 26551 17554 26560
rect 17604 26382 17632 28970
rect 17592 26376 17644 26382
rect 17592 26318 17644 26324
rect 17408 25696 17460 25702
rect 17408 25638 17460 25644
rect 17696 25226 17724 30330
rect 17868 30252 17920 30258
rect 17868 30194 17920 30200
rect 17880 29782 17908 30194
rect 17868 29776 17920 29782
rect 17868 29718 17920 29724
rect 17776 29572 17828 29578
rect 17776 29514 17828 29520
rect 17788 29170 17816 29514
rect 17776 29164 17828 29170
rect 17776 29106 17828 29112
rect 17788 28558 17816 29106
rect 17776 28552 17828 28558
rect 17776 28494 17828 28500
rect 17972 27849 18000 31146
rect 18052 31136 18104 31142
rect 18052 31078 18104 31084
rect 18144 31136 18196 31142
rect 18144 31078 18196 31084
rect 18064 30258 18092 31078
rect 18052 30252 18104 30258
rect 18052 30194 18104 30200
rect 18052 30048 18104 30054
rect 18052 29990 18104 29996
rect 18064 29594 18092 29990
rect 18156 29782 18184 31078
rect 18248 30122 18276 33200
rect 20456 31754 20484 33200
rect 19708 31748 19760 31754
rect 20456 31726 20760 31754
rect 19708 31690 19760 31696
rect 19720 31278 19748 31690
rect 20732 31346 20760 31726
rect 21364 31408 21416 31414
rect 21364 31350 21416 31356
rect 20444 31340 20496 31346
rect 20444 31282 20496 31288
rect 20536 31340 20588 31346
rect 20536 31282 20588 31288
rect 20720 31340 20772 31346
rect 20720 31282 20772 31288
rect 19708 31272 19760 31278
rect 18694 31240 18750 31249
rect 19708 31214 19760 31220
rect 18694 31175 18750 31184
rect 18315 31036 18623 31045
rect 18315 31034 18321 31036
rect 18377 31034 18401 31036
rect 18457 31034 18481 31036
rect 18537 31034 18561 31036
rect 18617 31034 18623 31036
rect 18377 30982 18379 31034
rect 18559 30982 18561 31034
rect 18315 30980 18321 30982
rect 18377 30980 18401 30982
rect 18457 30980 18481 30982
rect 18537 30980 18561 30982
rect 18617 30980 18623 30982
rect 18315 30971 18623 30980
rect 18236 30116 18288 30122
rect 18236 30058 18288 30064
rect 18315 29948 18623 29957
rect 18315 29946 18321 29948
rect 18377 29946 18401 29948
rect 18457 29946 18481 29948
rect 18537 29946 18561 29948
rect 18617 29946 18623 29948
rect 18377 29894 18379 29946
rect 18559 29894 18561 29946
rect 18315 29892 18321 29894
rect 18377 29892 18401 29894
rect 18457 29892 18481 29894
rect 18537 29892 18561 29894
rect 18617 29892 18623 29894
rect 18315 29883 18623 29892
rect 18708 29782 18736 31175
rect 19616 31136 19668 31142
rect 19616 31078 19668 31084
rect 18788 30864 18840 30870
rect 18788 30806 18840 30812
rect 18144 29776 18196 29782
rect 18696 29776 18748 29782
rect 18196 29724 18276 29730
rect 18144 29718 18276 29724
rect 18696 29718 18748 29724
rect 18156 29702 18276 29718
rect 18064 29566 18184 29594
rect 18052 29504 18104 29510
rect 18052 29446 18104 29452
rect 18064 29306 18092 29446
rect 18052 29300 18104 29306
rect 18052 29242 18104 29248
rect 18156 28801 18184 29566
rect 18142 28792 18198 28801
rect 18142 28727 18198 28736
rect 18156 28694 18184 28727
rect 18144 28688 18196 28694
rect 18144 28630 18196 28636
rect 17958 27840 18014 27849
rect 17958 27775 18014 27784
rect 18248 26586 18276 29702
rect 18696 29640 18748 29646
rect 18696 29582 18748 29588
rect 18315 28860 18623 28869
rect 18315 28858 18321 28860
rect 18377 28858 18401 28860
rect 18457 28858 18481 28860
rect 18537 28858 18561 28860
rect 18617 28858 18623 28860
rect 18377 28806 18379 28858
rect 18559 28806 18561 28858
rect 18315 28804 18321 28806
rect 18377 28804 18401 28806
rect 18457 28804 18481 28806
rect 18537 28804 18561 28806
rect 18617 28804 18623 28806
rect 18315 28795 18623 28804
rect 18708 28762 18736 29582
rect 18800 29034 18828 30806
rect 19260 30802 19564 30818
rect 19248 30796 19564 30802
rect 19300 30790 19564 30796
rect 19248 30738 19300 30744
rect 19536 30734 19564 30790
rect 19064 30728 19116 30734
rect 19064 30670 19116 30676
rect 19524 30728 19576 30734
rect 19524 30670 19576 30676
rect 18972 30048 19024 30054
rect 18972 29990 19024 29996
rect 18880 29640 18932 29646
rect 18984 29617 19012 29990
rect 18880 29582 18932 29588
rect 18970 29608 19026 29617
rect 18788 29028 18840 29034
rect 18788 28970 18840 28976
rect 18696 28756 18748 28762
rect 18696 28698 18748 28704
rect 18892 27878 18920 29582
rect 18970 29543 19026 29552
rect 19076 29345 19104 30670
rect 19628 30326 19656 31078
rect 19720 30666 19748 31214
rect 20168 31204 20220 31210
rect 20168 31146 20220 31152
rect 19892 31136 19944 31142
rect 19892 31078 19944 31084
rect 19800 30864 19852 30870
rect 19798 30832 19800 30841
rect 19852 30832 19854 30841
rect 19798 30767 19854 30776
rect 19708 30660 19760 30666
rect 19708 30602 19760 30608
rect 19904 30433 19932 31078
rect 20180 30734 20208 31146
rect 20456 30938 20484 31282
rect 20444 30932 20496 30938
rect 20444 30874 20496 30880
rect 20168 30728 20220 30734
rect 20168 30670 20220 30676
rect 20352 30728 20404 30734
rect 20352 30670 20404 30676
rect 20260 30592 20312 30598
rect 20260 30534 20312 30540
rect 19890 30424 19946 30433
rect 19890 30359 19946 30368
rect 19616 30320 19668 30326
rect 19616 30262 19668 30268
rect 19524 30252 19576 30258
rect 19524 30194 19576 30200
rect 19536 29578 19564 30194
rect 19628 30161 19656 30262
rect 19614 30152 19670 30161
rect 19614 30087 19670 30096
rect 20272 29850 20300 30534
rect 20260 29844 20312 29850
rect 20260 29786 20312 29792
rect 20364 29578 20392 30670
rect 20548 30666 20576 31282
rect 21376 30938 21404 31350
rect 21560 31346 21588 33200
rect 21788 31580 22096 31589
rect 21788 31578 21794 31580
rect 21850 31578 21874 31580
rect 21930 31578 21954 31580
rect 22010 31578 22034 31580
rect 22090 31578 22096 31580
rect 21850 31526 21852 31578
rect 22032 31526 22034 31578
rect 21788 31524 21794 31526
rect 21850 31524 21874 31526
rect 21930 31524 21954 31526
rect 22010 31524 22034 31526
rect 22090 31524 22096 31526
rect 21788 31515 22096 31524
rect 23768 31346 23796 33200
rect 24872 31346 24900 33200
rect 27080 31346 27108 33200
rect 27710 31920 27766 31929
rect 27710 31855 27766 31864
rect 21548 31340 21600 31346
rect 21548 31282 21600 31288
rect 23756 31340 23808 31346
rect 23756 31282 23808 31288
rect 24860 31340 24912 31346
rect 24860 31282 24912 31288
rect 27068 31340 27120 31346
rect 27068 31282 27120 31288
rect 25261 31036 25569 31045
rect 25261 31034 25267 31036
rect 25323 31034 25347 31036
rect 25403 31034 25427 31036
rect 25483 31034 25507 31036
rect 25563 31034 25569 31036
rect 25323 30982 25325 31034
rect 25505 30982 25507 31034
rect 25261 30980 25267 30982
rect 25323 30980 25347 30982
rect 25403 30980 25427 30982
rect 25483 30980 25507 30982
rect 25563 30980 25569 30982
rect 25261 30971 25569 30980
rect 27724 30938 27752 31855
rect 28184 31346 28212 33200
rect 28734 31580 29042 31589
rect 28734 31578 28740 31580
rect 28796 31578 28820 31580
rect 28876 31578 28900 31580
rect 28956 31578 28980 31580
rect 29036 31578 29042 31580
rect 28796 31526 28798 31578
rect 28978 31526 28980 31578
rect 28734 31524 28740 31526
rect 28796 31524 28820 31526
rect 28876 31524 28900 31526
rect 28956 31524 28980 31526
rect 29036 31524 29042 31526
rect 28734 31515 29042 31524
rect 28172 31340 28224 31346
rect 28172 31282 28224 31288
rect 28354 31240 28410 31249
rect 28354 31175 28410 31184
rect 28368 30938 28396 31175
rect 21364 30932 21416 30938
rect 21364 30874 21416 30880
rect 27712 30932 27764 30938
rect 27712 30874 27764 30880
rect 28356 30932 28408 30938
rect 28356 30874 28408 30880
rect 20536 30660 20588 30666
rect 20536 30602 20588 30608
rect 21788 30492 22096 30501
rect 21788 30490 21794 30492
rect 21850 30490 21874 30492
rect 21930 30490 21954 30492
rect 22010 30490 22034 30492
rect 22090 30490 22096 30492
rect 21850 30438 21852 30490
rect 22032 30438 22034 30490
rect 21788 30436 21794 30438
rect 21850 30436 21874 30438
rect 21930 30436 21954 30438
rect 22010 30436 22034 30438
rect 22090 30436 22096 30438
rect 21788 30427 22096 30436
rect 28734 30492 29042 30501
rect 28734 30490 28740 30492
rect 28796 30490 28820 30492
rect 28876 30490 28900 30492
rect 28956 30490 28980 30492
rect 29036 30490 29042 30492
rect 28796 30438 28798 30490
rect 28978 30438 28980 30490
rect 28734 30436 28740 30438
rect 28796 30436 28820 30438
rect 28876 30436 28900 30438
rect 28956 30436 28980 30438
rect 29036 30436 29042 30438
rect 28734 30427 29042 30436
rect 28356 30048 28408 30054
rect 28356 29990 28408 29996
rect 25261 29948 25569 29957
rect 25261 29946 25267 29948
rect 25323 29946 25347 29948
rect 25403 29946 25427 29948
rect 25483 29946 25507 29948
rect 25563 29946 25569 29948
rect 25323 29894 25325 29946
rect 25505 29894 25507 29946
rect 25261 29892 25267 29894
rect 25323 29892 25347 29894
rect 25403 29892 25427 29894
rect 25483 29892 25507 29894
rect 25563 29892 25569 29894
rect 25261 29883 25569 29892
rect 28368 29889 28396 29990
rect 28354 29880 28410 29889
rect 28354 29815 28410 29824
rect 28356 29640 28408 29646
rect 28356 29582 28408 29588
rect 19524 29572 19576 29578
rect 19524 29514 19576 29520
rect 20352 29572 20404 29578
rect 20352 29514 20404 29520
rect 21788 29404 22096 29413
rect 21788 29402 21794 29404
rect 21850 29402 21874 29404
rect 21930 29402 21954 29404
rect 22010 29402 22034 29404
rect 22090 29402 22096 29404
rect 21850 29350 21852 29402
rect 22032 29350 22034 29402
rect 21788 29348 21794 29350
rect 21850 29348 21874 29350
rect 21930 29348 21954 29350
rect 22010 29348 22034 29350
rect 22090 29348 22096 29350
rect 19062 29336 19118 29345
rect 21788 29339 22096 29348
rect 19062 29271 19118 29280
rect 28368 29209 28396 29582
rect 28734 29404 29042 29413
rect 28734 29402 28740 29404
rect 28796 29402 28820 29404
rect 28876 29402 28900 29404
rect 28956 29402 28980 29404
rect 29036 29402 29042 29404
rect 28796 29350 28798 29402
rect 28978 29350 28980 29402
rect 28734 29348 28740 29350
rect 28796 29348 28820 29350
rect 28876 29348 28900 29350
rect 28956 29348 28980 29350
rect 29036 29348 29042 29350
rect 28734 29339 29042 29348
rect 28354 29200 28410 29209
rect 28354 29135 28410 29144
rect 25261 28860 25569 28869
rect 25261 28858 25267 28860
rect 25323 28858 25347 28860
rect 25403 28858 25427 28860
rect 25483 28858 25507 28860
rect 25563 28858 25569 28860
rect 25323 28806 25325 28858
rect 25505 28806 25507 28858
rect 25261 28804 25267 28806
rect 25323 28804 25347 28806
rect 25403 28804 25427 28806
rect 25483 28804 25507 28806
rect 25563 28804 25569 28806
rect 25261 28795 25569 28804
rect 21788 28316 22096 28325
rect 21788 28314 21794 28316
rect 21850 28314 21874 28316
rect 21930 28314 21954 28316
rect 22010 28314 22034 28316
rect 22090 28314 22096 28316
rect 21850 28262 21852 28314
rect 22032 28262 22034 28314
rect 21788 28260 21794 28262
rect 21850 28260 21874 28262
rect 21930 28260 21954 28262
rect 22010 28260 22034 28262
rect 22090 28260 22096 28262
rect 21788 28251 22096 28260
rect 28734 28316 29042 28325
rect 28734 28314 28740 28316
rect 28796 28314 28820 28316
rect 28876 28314 28900 28316
rect 28956 28314 28980 28316
rect 29036 28314 29042 28316
rect 28796 28262 28798 28314
rect 28978 28262 28980 28314
rect 28734 28260 28740 28262
rect 28796 28260 28820 28262
rect 28876 28260 28900 28262
rect 28956 28260 28980 28262
rect 29036 28260 29042 28262
rect 28734 28251 29042 28260
rect 18880 27872 18932 27878
rect 28356 27872 28408 27878
rect 18880 27814 18932 27820
rect 28354 27840 28356 27849
rect 28408 27840 28410 27849
rect 18315 27772 18623 27781
rect 18315 27770 18321 27772
rect 18377 27770 18401 27772
rect 18457 27770 18481 27772
rect 18537 27770 18561 27772
rect 18617 27770 18623 27772
rect 18377 27718 18379 27770
rect 18559 27718 18561 27770
rect 18315 27716 18321 27718
rect 18377 27716 18401 27718
rect 18457 27716 18481 27718
rect 18537 27716 18561 27718
rect 18617 27716 18623 27718
rect 18315 27707 18623 27716
rect 25261 27772 25569 27781
rect 28354 27775 28410 27784
rect 25261 27770 25267 27772
rect 25323 27770 25347 27772
rect 25403 27770 25427 27772
rect 25483 27770 25507 27772
rect 25563 27770 25569 27772
rect 25323 27718 25325 27770
rect 25505 27718 25507 27770
rect 25261 27716 25267 27718
rect 25323 27716 25347 27718
rect 25403 27716 25427 27718
rect 25483 27716 25507 27718
rect 25563 27716 25569 27718
rect 25261 27707 25569 27716
rect 28356 27464 28408 27470
rect 28354 27432 28356 27441
rect 28408 27432 28410 27441
rect 28354 27367 28410 27376
rect 21788 27228 22096 27237
rect 21788 27226 21794 27228
rect 21850 27226 21874 27228
rect 21930 27226 21954 27228
rect 22010 27226 22034 27228
rect 22090 27226 22096 27228
rect 21850 27174 21852 27226
rect 22032 27174 22034 27226
rect 21788 27172 21794 27174
rect 21850 27172 21874 27174
rect 21930 27172 21954 27174
rect 22010 27172 22034 27174
rect 22090 27172 22096 27174
rect 21788 27163 22096 27172
rect 28734 27228 29042 27237
rect 28734 27226 28740 27228
rect 28796 27226 28820 27228
rect 28876 27226 28900 27228
rect 28956 27226 28980 27228
rect 29036 27226 29042 27228
rect 28796 27174 28798 27226
rect 28978 27174 28980 27226
rect 28734 27172 28740 27174
rect 28796 27172 28820 27174
rect 28876 27172 28900 27174
rect 28956 27172 28980 27174
rect 29036 27172 29042 27174
rect 28734 27163 29042 27172
rect 18315 26684 18623 26693
rect 18315 26682 18321 26684
rect 18377 26682 18401 26684
rect 18457 26682 18481 26684
rect 18537 26682 18561 26684
rect 18617 26682 18623 26684
rect 18377 26630 18379 26682
rect 18559 26630 18561 26682
rect 18315 26628 18321 26630
rect 18377 26628 18401 26630
rect 18457 26628 18481 26630
rect 18537 26628 18561 26630
rect 18617 26628 18623 26630
rect 18315 26619 18623 26628
rect 25261 26684 25569 26693
rect 25261 26682 25267 26684
rect 25323 26682 25347 26684
rect 25403 26682 25427 26684
rect 25483 26682 25507 26684
rect 25563 26682 25569 26684
rect 25323 26630 25325 26682
rect 25505 26630 25507 26682
rect 25261 26628 25267 26630
rect 25323 26628 25347 26630
rect 25403 26628 25427 26630
rect 25483 26628 25507 26630
rect 25563 26628 25569 26630
rect 25261 26619 25569 26628
rect 18236 26580 18288 26586
rect 18236 26522 18288 26528
rect 21788 26140 22096 26149
rect 21788 26138 21794 26140
rect 21850 26138 21874 26140
rect 21930 26138 21954 26140
rect 22010 26138 22034 26140
rect 22090 26138 22096 26140
rect 21850 26086 21852 26138
rect 22032 26086 22034 26138
rect 21788 26084 21794 26086
rect 21850 26084 21874 26086
rect 21930 26084 21954 26086
rect 22010 26084 22034 26086
rect 22090 26084 22096 26086
rect 21788 26075 22096 26084
rect 28734 26140 29042 26149
rect 28734 26138 28740 26140
rect 28796 26138 28820 26140
rect 28876 26138 28900 26140
rect 28956 26138 28980 26140
rect 29036 26138 29042 26140
rect 28796 26086 28798 26138
rect 28978 26086 28980 26138
rect 28734 26084 28740 26086
rect 28796 26084 28820 26086
rect 28876 26084 28900 26086
rect 28956 26084 28980 26086
rect 29036 26084 29042 26086
rect 28734 26075 29042 26084
rect 28354 25800 28410 25809
rect 28354 25735 28356 25744
rect 28408 25735 28410 25744
rect 28356 25706 28408 25712
rect 18315 25596 18623 25605
rect 18315 25594 18321 25596
rect 18377 25594 18401 25596
rect 18457 25594 18481 25596
rect 18537 25594 18561 25596
rect 18617 25594 18623 25596
rect 18377 25542 18379 25594
rect 18559 25542 18561 25594
rect 18315 25540 18321 25542
rect 18377 25540 18401 25542
rect 18457 25540 18481 25542
rect 18537 25540 18561 25542
rect 18617 25540 18623 25542
rect 18315 25531 18623 25540
rect 25261 25596 25569 25605
rect 25261 25594 25267 25596
rect 25323 25594 25347 25596
rect 25403 25594 25427 25596
rect 25483 25594 25507 25596
rect 25563 25594 25569 25596
rect 25323 25542 25325 25594
rect 25505 25542 25507 25594
rect 25261 25540 25267 25542
rect 25323 25540 25347 25542
rect 25403 25540 25427 25542
rect 25483 25540 25507 25542
rect 25563 25540 25569 25542
rect 25261 25531 25569 25540
rect 28356 25424 28408 25430
rect 28354 25392 28356 25401
rect 28408 25392 28410 25401
rect 28354 25327 28410 25336
rect 17684 25220 17736 25226
rect 17684 25162 17736 25168
rect 21788 25052 22096 25061
rect 21788 25050 21794 25052
rect 21850 25050 21874 25052
rect 21930 25050 21954 25052
rect 22010 25050 22034 25052
rect 22090 25050 22096 25052
rect 21850 24998 21852 25050
rect 22032 24998 22034 25050
rect 21788 24996 21794 24998
rect 21850 24996 21874 24998
rect 21930 24996 21954 24998
rect 22010 24996 22034 24998
rect 22090 24996 22096 24998
rect 21788 24987 22096 24996
rect 28734 25052 29042 25061
rect 28734 25050 28740 25052
rect 28796 25050 28820 25052
rect 28876 25050 28900 25052
rect 28956 25050 28980 25052
rect 29036 25050 29042 25052
rect 28796 24998 28798 25050
rect 28978 24998 28980 25050
rect 28734 24996 28740 24998
rect 28796 24996 28820 24998
rect 28876 24996 28900 24998
rect 28956 24996 28980 24998
rect 29036 24996 29042 24998
rect 28734 24987 29042 24996
rect 18315 24508 18623 24517
rect 18315 24506 18321 24508
rect 18377 24506 18401 24508
rect 18457 24506 18481 24508
rect 18537 24506 18561 24508
rect 18617 24506 18623 24508
rect 18377 24454 18379 24506
rect 18559 24454 18561 24506
rect 18315 24452 18321 24454
rect 18377 24452 18401 24454
rect 18457 24452 18481 24454
rect 18537 24452 18561 24454
rect 18617 24452 18623 24454
rect 18315 24443 18623 24452
rect 25261 24508 25569 24517
rect 25261 24506 25267 24508
rect 25323 24506 25347 24508
rect 25403 24506 25427 24508
rect 25483 24506 25507 24508
rect 25563 24506 25569 24508
rect 25323 24454 25325 24506
rect 25505 24454 25507 24506
rect 25261 24452 25267 24454
rect 25323 24452 25347 24454
rect 25403 24452 25427 24454
rect 25483 24452 25507 24454
rect 25563 24452 25569 24454
rect 25261 24443 25569 24452
rect 28356 24200 28408 24206
rect 28356 24142 28408 24148
rect 21788 23964 22096 23973
rect 21788 23962 21794 23964
rect 21850 23962 21874 23964
rect 21930 23962 21954 23964
rect 22010 23962 22034 23964
rect 22090 23962 22096 23964
rect 21850 23910 21852 23962
rect 22032 23910 22034 23962
rect 21788 23908 21794 23910
rect 21850 23908 21874 23910
rect 21930 23908 21954 23910
rect 22010 23908 22034 23910
rect 22090 23908 22096 23910
rect 21788 23899 22096 23908
rect 28368 23769 28396 24142
rect 28734 23964 29042 23973
rect 28734 23962 28740 23964
rect 28796 23962 28820 23964
rect 28876 23962 28900 23964
rect 28956 23962 28980 23964
rect 29036 23962 29042 23964
rect 28796 23910 28798 23962
rect 28978 23910 28980 23962
rect 28734 23908 28740 23910
rect 28796 23908 28820 23910
rect 28876 23908 28900 23910
rect 28956 23908 28980 23910
rect 29036 23908 29042 23910
rect 28734 23899 29042 23908
rect 28354 23760 28410 23769
rect 28354 23695 28410 23704
rect 18315 23420 18623 23429
rect 18315 23418 18321 23420
rect 18377 23418 18401 23420
rect 18457 23418 18481 23420
rect 18537 23418 18561 23420
rect 18617 23418 18623 23420
rect 18377 23366 18379 23418
rect 18559 23366 18561 23418
rect 18315 23364 18321 23366
rect 18377 23364 18401 23366
rect 18457 23364 18481 23366
rect 18537 23364 18561 23366
rect 18617 23364 18623 23366
rect 18315 23355 18623 23364
rect 25261 23420 25569 23429
rect 25261 23418 25267 23420
rect 25323 23418 25347 23420
rect 25403 23418 25427 23420
rect 25483 23418 25507 23420
rect 25563 23418 25569 23420
rect 25323 23366 25325 23418
rect 25505 23366 25507 23418
rect 25261 23364 25267 23366
rect 25323 23364 25347 23366
rect 25403 23364 25427 23366
rect 25483 23364 25507 23366
rect 25563 23364 25569 23366
rect 25261 23355 25569 23364
rect 28356 23112 28408 23118
rect 28354 23080 28356 23089
rect 28408 23080 28410 23089
rect 28354 23015 28410 23024
rect 21788 22876 22096 22885
rect 21788 22874 21794 22876
rect 21850 22874 21874 22876
rect 21930 22874 21954 22876
rect 22010 22874 22034 22876
rect 22090 22874 22096 22876
rect 21850 22822 21852 22874
rect 22032 22822 22034 22874
rect 21788 22820 21794 22822
rect 21850 22820 21874 22822
rect 21930 22820 21954 22822
rect 22010 22820 22034 22822
rect 22090 22820 22096 22822
rect 21788 22811 22096 22820
rect 28734 22876 29042 22885
rect 28734 22874 28740 22876
rect 28796 22874 28820 22876
rect 28876 22874 28900 22876
rect 28956 22874 28980 22876
rect 29036 22874 29042 22876
rect 28796 22822 28798 22874
rect 28978 22822 28980 22874
rect 28734 22820 28740 22822
rect 28796 22820 28820 22822
rect 28876 22820 28900 22822
rect 28956 22820 28980 22822
rect 29036 22820 29042 22822
rect 28734 22811 29042 22820
rect 18315 22332 18623 22341
rect 18315 22330 18321 22332
rect 18377 22330 18401 22332
rect 18457 22330 18481 22332
rect 18537 22330 18561 22332
rect 18617 22330 18623 22332
rect 18377 22278 18379 22330
rect 18559 22278 18561 22330
rect 18315 22276 18321 22278
rect 18377 22276 18401 22278
rect 18457 22276 18481 22278
rect 18537 22276 18561 22278
rect 18617 22276 18623 22278
rect 18315 22267 18623 22276
rect 25261 22332 25569 22341
rect 25261 22330 25267 22332
rect 25323 22330 25347 22332
rect 25403 22330 25427 22332
rect 25483 22330 25507 22332
rect 25563 22330 25569 22332
rect 25323 22278 25325 22330
rect 25505 22278 25507 22330
rect 25261 22276 25267 22278
rect 25323 22276 25347 22278
rect 25403 22276 25427 22278
rect 25483 22276 25507 22278
rect 25563 22276 25569 22278
rect 25261 22267 25569 22276
rect 28356 22024 28408 22030
rect 28354 21992 28356 22001
rect 28408 21992 28410 22001
rect 28354 21927 28410 21936
rect 21788 21788 22096 21797
rect 21788 21786 21794 21788
rect 21850 21786 21874 21788
rect 21930 21786 21954 21788
rect 22010 21786 22034 21788
rect 22090 21786 22096 21788
rect 21850 21734 21852 21786
rect 22032 21734 22034 21786
rect 21788 21732 21794 21734
rect 21850 21732 21874 21734
rect 21930 21732 21954 21734
rect 22010 21732 22034 21734
rect 22090 21732 22096 21734
rect 21788 21723 22096 21732
rect 28734 21788 29042 21797
rect 28734 21786 28740 21788
rect 28796 21786 28820 21788
rect 28876 21786 28900 21788
rect 28956 21786 28980 21788
rect 29036 21786 29042 21788
rect 28796 21734 28798 21786
rect 28978 21734 28980 21786
rect 28734 21732 28740 21734
rect 28796 21732 28820 21734
rect 28876 21732 28900 21734
rect 28956 21732 28980 21734
rect 29036 21732 29042 21734
rect 28734 21723 29042 21732
rect 28356 21344 28408 21350
rect 28356 21286 28408 21292
rect 18315 21244 18623 21253
rect 18315 21242 18321 21244
rect 18377 21242 18401 21244
rect 18457 21242 18481 21244
rect 18537 21242 18561 21244
rect 18617 21242 18623 21244
rect 18377 21190 18379 21242
rect 18559 21190 18561 21242
rect 18315 21188 18321 21190
rect 18377 21188 18401 21190
rect 18457 21188 18481 21190
rect 18537 21188 18561 21190
rect 18617 21188 18623 21190
rect 18315 21179 18623 21188
rect 25261 21244 25569 21253
rect 25261 21242 25267 21244
rect 25323 21242 25347 21244
rect 25403 21242 25427 21244
rect 25483 21242 25507 21244
rect 25563 21242 25569 21244
rect 25323 21190 25325 21242
rect 25505 21190 25507 21242
rect 25261 21188 25267 21190
rect 25323 21188 25347 21190
rect 25403 21188 25427 21190
rect 25483 21188 25507 21190
rect 25563 21188 25569 21190
rect 25261 21179 25569 21188
rect 28368 21049 28396 21286
rect 28354 21040 28410 21049
rect 28354 20975 28410 20984
rect 21788 20700 22096 20709
rect 21788 20698 21794 20700
rect 21850 20698 21874 20700
rect 21930 20698 21954 20700
rect 22010 20698 22034 20700
rect 22090 20698 22096 20700
rect 21850 20646 21852 20698
rect 22032 20646 22034 20698
rect 21788 20644 21794 20646
rect 21850 20644 21874 20646
rect 21930 20644 21954 20646
rect 22010 20644 22034 20646
rect 22090 20644 22096 20646
rect 21788 20635 22096 20644
rect 28734 20700 29042 20709
rect 28734 20698 28740 20700
rect 28796 20698 28820 20700
rect 28876 20698 28900 20700
rect 28956 20698 28980 20700
rect 29036 20698 29042 20700
rect 28796 20646 28798 20698
rect 28978 20646 28980 20698
rect 28734 20644 28740 20646
rect 28796 20644 28820 20646
rect 28876 20644 28900 20646
rect 28956 20644 28980 20646
rect 29036 20644 29042 20646
rect 28734 20635 29042 20644
rect 18315 20156 18623 20165
rect 18315 20154 18321 20156
rect 18377 20154 18401 20156
rect 18457 20154 18481 20156
rect 18537 20154 18561 20156
rect 18617 20154 18623 20156
rect 18377 20102 18379 20154
rect 18559 20102 18561 20154
rect 18315 20100 18321 20102
rect 18377 20100 18401 20102
rect 18457 20100 18481 20102
rect 18537 20100 18561 20102
rect 18617 20100 18623 20102
rect 18315 20091 18623 20100
rect 25261 20156 25569 20165
rect 25261 20154 25267 20156
rect 25323 20154 25347 20156
rect 25403 20154 25427 20156
rect 25483 20154 25507 20156
rect 25563 20154 25569 20156
rect 25323 20102 25325 20154
rect 25505 20102 25507 20154
rect 25261 20100 25267 20102
rect 25323 20100 25347 20102
rect 25403 20100 25427 20102
rect 25483 20100 25507 20102
rect 25563 20100 25569 20102
rect 25261 20091 25569 20100
rect 28356 19984 28408 19990
rect 28354 19952 28356 19961
rect 28408 19952 28410 19961
rect 28354 19887 28410 19896
rect 21788 19612 22096 19621
rect 21788 19610 21794 19612
rect 21850 19610 21874 19612
rect 21930 19610 21954 19612
rect 22010 19610 22034 19612
rect 22090 19610 22096 19612
rect 21850 19558 21852 19610
rect 22032 19558 22034 19610
rect 21788 19556 21794 19558
rect 21850 19556 21874 19558
rect 21930 19556 21954 19558
rect 22010 19556 22034 19558
rect 22090 19556 22096 19558
rect 21788 19547 22096 19556
rect 28734 19612 29042 19621
rect 28734 19610 28740 19612
rect 28796 19610 28820 19612
rect 28876 19610 28900 19612
rect 28956 19610 28980 19612
rect 29036 19610 29042 19612
rect 28796 19558 28798 19610
rect 28978 19558 28980 19610
rect 28734 19556 28740 19558
rect 28796 19556 28820 19558
rect 28876 19556 28900 19558
rect 28956 19556 28980 19558
rect 29036 19556 29042 19558
rect 28734 19547 29042 19556
rect 28356 19168 28408 19174
rect 28356 19110 28408 19116
rect 18315 19068 18623 19077
rect 18315 19066 18321 19068
rect 18377 19066 18401 19068
rect 18457 19066 18481 19068
rect 18537 19066 18561 19068
rect 18617 19066 18623 19068
rect 18377 19014 18379 19066
rect 18559 19014 18561 19066
rect 18315 19012 18321 19014
rect 18377 19012 18401 19014
rect 18457 19012 18481 19014
rect 18537 19012 18561 19014
rect 18617 19012 18623 19014
rect 18315 19003 18623 19012
rect 25261 19068 25569 19077
rect 25261 19066 25267 19068
rect 25323 19066 25347 19068
rect 25403 19066 25427 19068
rect 25483 19066 25507 19068
rect 25563 19066 25569 19068
rect 25323 19014 25325 19066
rect 25505 19014 25507 19066
rect 25261 19012 25267 19014
rect 25323 19012 25347 19014
rect 25403 19012 25427 19014
rect 25483 19012 25507 19014
rect 25563 19012 25569 19014
rect 25261 19003 25569 19012
rect 28368 19009 28396 19110
rect 28354 19000 28410 19009
rect 28354 18935 28410 18944
rect 21788 18524 22096 18533
rect 21788 18522 21794 18524
rect 21850 18522 21874 18524
rect 21930 18522 21954 18524
rect 22010 18522 22034 18524
rect 22090 18522 22096 18524
rect 21850 18470 21852 18522
rect 22032 18470 22034 18522
rect 21788 18468 21794 18470
rect 21850 18468 21874 18470
rect 21930 18468 21954 18470
rect 22010 18468 22034 18470
rect 22090 18468 22096 18470
rect 21788 18459 22096 18468
rect 28734 18524 29042 18533
rect 28734 18522 28740 18524
rect 28796 18522 28820 18524
rect 28876 18522 28900 18524
rect 28956 18522 28980 18524
rect 29036 18522 29042 18524
rect 28796 18470 28798 18522
rect 28978 18470 28980 18522
rect 28734 18468 28740 18470
rect 28796 18468 28820 18470
rect 28876 18468 28900 18470
rect 28956 18468 28980 18470
rect 29036 18468 29042 18470
rect 28734 18459 29042 18468
rect 18315 17980 18623 17989
rect 18315 17978 18321 17980
rect 18377 17978 18401 17980
rect 18457 17978 18481 17980
rect 18537 17978 18561 17980
rect 18617 17978 18623 17980
rect 18377 17926 18379 17978
rect 18559 17926 18561 17978
rect 18315 17924 18321 17926
rect 18377 17924 18401 17926
rect 18457 17924 18481 17926
rect 18537 17924 18561 17926
rect 18617 17924 18623 17926
rect 18315 17915 18623 17924
rect 25261 17980 25569 17989
rect 25261 17978 25267 17980
rect 25323 17978 25347 17980
rect 25403 17978 25427 17980
rect 25483 17978 25507 17980
rect 25563 17978 25569 17980
rect 25323 17926 25325 17978
rect 25505 17926 25507 17978
rect 25261 17924 25267 17926
rect 25323 17924 25347 17926
rect 25403 17924 25427 17926
rect 25483 17924 25507 17926
rect 25563 17924 25569 17926
rect 25261 17915 25569 17924
rect 28356 17672 28408 17678
rect 28354 17640 28356 17649
rect 28408 17640 28410 17649
rect 28354 17575 28410 17584
rect 21788 17436 22096 17445
rect 21788 17434 21794 17436
rect 21850 17434 21874 17436
rect 21930 17434 21954 17436
rect 22010 17434 22034 17436
rect 22090 17434 22096 17436
rect 21850 17382 21852 17434
rect 22032 17382 22034 17434
rect 21788 17380 21794 17382
rect 21850 17380 21874 17382
rect 21930 17380 21954 17382
rect 22010 17380 22034 17382
rect 22090 17380 22096 17382
rect 21788 17371 22096 17380
rect 28734 17436 29042 17445
rect 28734 17434 28740 17436
rect 28796 17434 28820 17436
rect 28876 17434 28900 17436
rect 28956 17434 28980 17436
rect 29036 17434 29042 17436
rect 28796 17382 28798 17434
rect 28978 17382 28980 17434
rect 28734 17380 28740 17382
rect 28796 17380 28820 17382
rect 28876 17380 28900 17382
rect 28956 17380 28980 17382
rect 29036 17380 29042 17382
rect 28734 17371 29042 17380
rect 28356 16992 28408 16998
rect 28354 16960 28356 16969
rect 28408 16960 28410 16969
rect 18315 16892 18623 16901
rect 18315 16890 18321 16892
rect 18377 16890 18401 16892
rect 18457 16890 18481 16892
rect 18537 16890 18561 16892
rect 18617 16890 18623 16892
rect 18377 16838 18379 16890
rect 18559 16838 18561 16890
rect 18315 16836 18321 16838
rect 18377 16836 18401 16838
rect 18457 16836 18481 16838
rect 18537 16836 18561 16838
rect 18617 16836 18623 16838
rect 18315 16827 18623 16836
rect 25261 16892 25569 16901
rect 28354 16895 28410 16904
rect 25261 16890 25267 16892
rect 25323 16890 25347 16892
rect 25403 16890 25427 16892
rect 25483 16890 25507 16892
rect 25563 16890 25569 16892
rect 25323 16838 25325 16890
rect 25505 16838 25507 16890
rect 25261 16836 25267 16838
rect 25323 16836 25347 16838
rect 25403 16836 25427 16838
rect 25483 16836 25507 16838
rect 25563 16836 25569 16838
rect 25261 16827 25569 16836
rect 21788 16348 22096 16357
rect 21788 16346 21794 16348
rect 21850 16346 21874 16348
rect 21930 16346 21954 16348
rect 22010 16346 22034 16348
rect 22090 16346 22096 16348
rect 21850 16294 21852 16346
rect 22032 16294 22034 16346
rect 21788 16292 21794 16294
rect 21850 16292 21874 16294
rect 21930 16292 21954 16294
rect 22010 16292 22034 16294
rect 22090 16292 22096 16294
rect 21788 16283 22096 16292
rect 28734 16348 29042 16357
rect 28734 16346 28740 16348
rect 28796 16346 28820 16348
rect 28876 16346 28900 16348
rect 28956 16346 28980 16348
rect 29036 16346 29042 16348
rect 28796 16294 28798 16346
rect 28978 16294 28980 16346
rect 28734 16292 28740 16294
rect 28796 16292 28820 16294
rect 28876 16292 28900 16294
rect 28956 16292 28980 16294
rect 29036 16292 29042 16294
rect 28734 16283 29042 16292
rect 28356 15904 28408 15910
rect 28356 15846 28408 15852
rect 18315 15804 18623 15813
rect 18315 15802 18321 15804
rect 18377 15802 18401 15804
rect 18457 15802 18481 15804
rect 18537 15802 18561 15804
rect 18617 15802 18623 15804
rect 18377 15750 18379 15802
rect 18559 15750 18561 15802
rect 18315 15748 18321 15750
rect 18377 15748 18401 15750
rect 18457 15748 18481 15750
rect 18537 15748 18561 15750
rect 18617 15748 18623 15750
rect 18315 15739 18623 15748
rect 25261 15804 25569 15813
rect 25261 15802 25267 15804
rect 25323 15802 25347 15804
rect 25403 15802 25427 15804
rect 25483 15802 25507 15804
rect 25563 15802 25569 15804
rect 25323 15750 25325 15802
rect 25505 15750 25507 15802
rect 25261 15748 25267 15750
rect 25323 15748 25347 15750
rect 25403 15748 25427 15750
rect 25483 15748 25507 15750
rect 25563 15748 25569 15750
rect 25261 15739 25569 15748
rect 28368 15609 28396 15846
rect 28354 15600 28410 15609
rect 28354 15535 28410 15544
rect 21788 15260 22096 15269
rect 21788 15258 21794 15260
rect 21850 15258 21874 15260
rect 21930 15258 21954 15260
rect 22010 15258 22034 15260
rect 22090 15258 22096 15260
rect 21850 15206 21852 15258
rect 22032 15206 22034 15258
rect 21788 15204 21794 15206
rect 21850 15204 21874 15206
rect 21930 15204 21954 15206
rect 22010 15204 22034 15206
rect 22090 15204 22096 15206
rect 21788 15195 22096 15204
rect 28734 15260 29042 15269
rect 28734 15258 28740 15260
rect 28796 15258 28820 15260
rect 28876 15258 28900 15260
rect 28956 15258 28980 15260
rect 29036 15258 29042 15260
rect 28796 15206 28798 15258
rect 28978 15206 28980 15258
rect 28734 15204 28740 15206
rect 28796 15204 28820 15206
rect 28876 15204 28900 15206
rect 28956 15204 28980 15206
rect 29036 15204 29042 15206
rect 28734 15195 29042 15204
rect 28354 14920 28410 14929
rect 28354 14855 28356 14864
rect 28408 14855 28410 14864
rect 28356 14826 28408 14832
rect 18315 14716 18623 14725
rect 18315 14714 18321 14716
rect 18377 14714 18401 14716
rect 18457 14714 18481 14716
rect 18537 14714 18561 14716
rect 18617 14714 18623 14716
rect 18377 14662 18379 14714
rect 18559 14662 18561 14714
rect 18315 14660 18321 14662
rect 18377 14660 18401 14662
rect 18457 14660 18481 14662
rect 18537 14660 18561 14662
rect 18617 14660 18623 14662
rect 18315 14651 18623 14660
rect 25261 14716 25569 14725
rect 25261 14714 25267 14716
rect 25323 14714 25347 14716
rect 25403 14714 25427 14716
rect 25483 14714 25507 14716
rect 25563 14714 25569 14716
rect 25323 14662 25325 14714
rect 25505 14662 25507 14714
rect 25261 14660 25267 14662
rect 25323 14660 25347 14662
rect 25403 14660 25427 14662
rect 25483 14660 25507 14662
rect 25563 14660 25569 14662
rect 25261 14651 25569 14660
rect 21788 14172 22096 14181
rect 21788 14170 21794 14172
rect 21850 14170 21874 14172
rect 21930 14170 21954 14172
rect 22010 14170 22034 14172
rect 22090 14170 22096 14172
rect 21850 14118 21852 14170
rect 22032 14118 22034 14170
rect 21788 14116 21794 14118
rect 21850 14116 21874 14118
rect 21930 14116 21954 14118
rect 22010 14116 22034 14118
rect 22090 14116 22096 14118
rect 21788 14107 22096 14116
rect 28734 14172 29042 14181
rect 28734 14170 28740 14172
rect 28796 14170 28820 14172
rect 28876 14170 28900 14172
rect 28956 14170 28980 14172
rect 29036 14170 29042 14172
rect 28796 14118 28798 14170
rect 28978 14118 28980 14170
rect 28734 14116 28740 14118
rect 28796 14116 28820 14118
rect 28876 14116 28900 14118
rect 28956 14116 28980 14118
rect 29036 14116 29042 14118
rect 28734 14107 29042 14116
rect 28356 13728 28408 13734
rect 28356 13670 28408 13676
rect 18315 13628 18623 13637
rect 18315 13626 18321 13628
rect 18377 13626 18401 13628
rect 18457 13626 18481 13628
rect 18537 13626 18561 13628
rect 18617 13626 18623 13628
rect 18377 13574 18379 13626
rect 18559 13574 18561 13626
rect 18315 13572 18321 13574
rect 18377 13572 18401 13574
rect 18457 13572 18481 13574
rect 18537 13572 18561 13574
rect 18617 13572 18623 13574
rect 18315 13563 18623 13572
rect 25261 13628 25569 13637
rect 25261 13626 25267 13628
rect 25323 13626 25347 13628
rect 25403 13626 25427 13628
rect 25483 13626 25507 13628
rect 25563 13626 25569 13628
rect 25323 13574 25325 13626
rect 25505 13574 25507 13626
rect 25261 13572 25267 13574
rect 25323 13572 25347 13574
rect 25403 13572 25427 13574
rect 25483 13572 25507 13574
rect 25563 13572 25569 13574
rect 25261 13563 25569 13572
rect 28368 13569 28396 13670
rect 28354 13560 28410 13569
rect 28354 13495 28410 13504
rect 28356 13320 28408 13326
rect 28356 13262 28408 13268
rect 21788 13084 22096 13093
rect 21788 13082 21794 13084
rect 21850 13082 21874 13084
rect 21930 13082 21954 13084
rect 22010 13082 22034 13084
rect 22090 13082 22096 13084
rect 21850 13030 21852 13082
rect 22032 13030 22034 13082
rect 21788 13028 21794 13030
rect 21850 13028 21874 13030
rect 21930 13028 21954 13030
rect 22010 13028 22034 13030
rect 22090 13028 22096 13030
rect 21788 13019 22096 13028
rect 28368 12889 28396 13262
rect 28734 13084 29042 13093
rect 28734 13082 28740 13084
rect 28796 13082 28820 13084
rect 28876 13082 28900 13084
rect 28956 13082 28980 13084
rect 29036 13082 29042 13084
rect 28796 13030 28798 13082
rect 28978 13030 28980 13082
rect 28734 13028 28740 13030
rect 28796 13028 28820 13030
rect 28876 13028 28900 13030
rect 28956 13028 28980 13030
rect 29036 13028 29042 13030
rect 28734 13019 29042 13028
rect 28354 12880 28410 12889
rect 28354 12815 28410 12824
rect 18315 12540 18623 12549
rect 18315 12538 18321 12540
rect 18377 12538 18401 12540
rect 18457 12538 18481 12540
rect 18537 12538 18561 12540
rect 18617 12538 18623 12540
rect 18377 12486 18379 12538
rect 18559 12486 18561 12538
rect 18315 12484 18321 12486
rect 18377 12484 18401 12486
rect 18457 12484 18481 12486
rect 18537 12484 18561 12486
rect 18617 12484 18623 12486
rect 18315 12475 18623 12484
rect 25261 12540 25569 12549
rect 25261 12538 25267 12540
rect 25323 12538 25347 12540
rect 25403 12538 25427 12540
rect 25483 12538 25507 12540
rect 25563 12538 25569 12540
rect 25323 12486 25325 12538
rect 25505 12486 25507 12538
rect 25261 12484 25267 12486
rect 25323 12484 25347 12486
rect 25403 12484 25427 12486
rect 25483 12484 25507 12486
rect 25563 12484 25569 12486
rect 25261 12475 25569 12484
rect 21788 11996 22096 12005
rect 21788 11994 21794 11996
rect 21850 11994 21874 11996
rect 21930 11994 21954 11996
rect 22010 11994 22034 11996
rect 22090 11994 22096 11996
rect 21850 11942 21852 11994
rect 22032 11942 22034 11994
rect 21788 11940 21794 11942
rect 21850 11940 21874 11942
rect 21930 11940 21954 11942
rect 22010 11940 22034 11942
rect 22090 11940 22096 11942
rect 21788 11931 22096 11940
rect 28734 11996 29042 12005
rect 28734 11994 28740 11996
rect 28796 11994 28820 11996
rect 28876 11994 28900 11996
rect 28956 11994 28980 11996
rect 29036 11994 29042 11996
rect 28796 11942 28798 11994
rect 28978 11942 28980 11994
rect 28734 11940 28740 11942
rect 28796 11940 28820 11942
rect 28876 11940 28900 11942
rect 28956 11940 28980 11942
rect 29036 11940 29042 11942
rect 28734 11931 29042 11940
rect 28356 11552 28408 11558
rect 28354 11520 28356 11529
rect 28408 11520 28410 11529
rect 18315 11452 18623 11461
rect 18315 11450 18321 11452
rect 18377 11450 18401 11452
rect 18457 11450 18481 11452
rect 18537 11450 18561 11452
rect 18617 11450 18623 11452
rect 18377 11398 18379 11450
rect 18559 11398 18561 11450
rect 18315 11396 18321 11398
rect 18377 11396 18401 11398
rect 18457 11396 18481 11398
rect 18537 11396 18561 11398
rect 18617 11396 18623 11398
rect 18315 11387 18623 11396
rect 25261 11452 25569 11461
rect 28354 11455 28410 11464
rect 25261 11450 25267 11452
rect 25323 11450 25347 11452
rect 25403 11450 25427 11452
rect 25483 11450 25507 11452
rect 25563 11450 25569 11452
rect 25323 11398 25325 11450
rect 25505 11398 25507 11450
rect 25261 11396 25267 11398
rect 25323 11396 25347 11398
rect 25403 11396 25427 11398
rect 25483 11396 25507 11398
rect 25563 11396 25569 11398
rect 25261 11387 25569 11396
rect 28356 11144 28408 11150
rect 28354 11112 28356 11121
rect 28408 11112 28410 11121
rect 28354 11047 28410 11056
rect 21788 10908 22096 10917
rect 21788 10906 21794 10908
rect 21850 10906 21874 10908
rect 21930 10906 21954 10908
rect 22010 10906 22034 10908
rect 22090 10906 22096 10908
rect 21850 10854 21852 10906
rect 22032 10854 22034 10906
rect 21788 10852 21794 10854
rect 21850 10852 21874 10854
rect 21930 10852 21954 10854
rect 22010 10852 22034 10854
rect 22090 10852 22096 10854
rect 21788 10843 22096 10852
rect 28734 10908 29042 10917
rect 28734 10906 28740 10908
rect 28796 10906 28820 10908
rect 28876 10906 28900 10908
rect 28956 10906 28980 10908
rect 29036 10906 29042 10908
rect 28796 10854 28798 10906
rect 28978 10854 28980 10906
rect 28734 10852 28740 10854
rect 28796 10852 28820 10854
rect 28876 10852 28900 10854
rect 28956 10852 28980 10854
rect 29036 10852 29042 10854
rect 28734 10843 29042 10852
rect 18315 10364 18623 10373
rect 18315 10362 18321 10364
rect 18377 10362 18401 10364
rect 18457 10362 18481 10364
rect 18537 10362 18561 10364
rect 18617 10362 18623 10364
rect 18377 10310 18379 10362
rect 18559 10310 18561 10362
rect 18315 10308 18321 10310
rect 18377 10308 18401 10310
rect 18457 10308 18481 10310
rect 18537 10308 18561 10310
rect 18617 10308 18623 10310
rect 18315 10299 18623 10308
rect 25261 10364 25569 10373
rect 25261 10362 25267 10364
rect 25323 10362 25347 10364
rect 25403 10362 25427 10364
rect 25483 10362 25507 10364
rect 25563 10362 25569 10364
rect 25323 10310 25325 10362
rect 25505 10310 25507 10362
rect 25261 10308 25267 10310
rect 25323 10308 25347 10310
rect 25403 10308 25427 10310
rect 25483 10308 25507 10310
rect 25563 10308 25569 10310
rect 25261 10299 25569 10308
rect 21788 9820 22096 9829
rect 21788 9818 21794 9820
rect 21850 9818 21874 9820
rect 21930 9818 21954 9820
rect 22010 9818 22034 9820
rect 22090 9818 22096 9820
rect 21850 9766 21852 9818
rect 22032 9766 22034 9818
rect 21788 9764 21794 9766
rect 21850 9764 21874 9766
rect 21930 9764 21954 9766
rect 22010 9764 22034 9766
rect 22090 9764 22096 9766
rect 21788 9755 22096 9764
rect 28734 9820 29042 9829
rect 28734 9818 28740 9820
rect 28796 9818 28820 9820
rect 28876 9818 28900 9820
rect 28956 9818 28980 9820
rect 29036 9818 29042 9820
rect 28796 9766 28798 9818
rect 28978 9766 28980 9818
rect 28734 9764 28740 9766
rect 28796 9764 28820 9766
rect 28876 9764 28900 9766
rect 28956 9764 28980 9766
rect 29036 9764 29042 9766
rect 28734 9755 29042 9764
rect 28354 9480 28410 9489
rect 28354 9415 28356 9424
rect 28408 9415 28410 9424
rect 28356 9386 28408 9392
rect 18315 9276 18623 9285
rect 18315 9274 18321 9276
rect 18377 9274 18401 9276
rect 18457 9274 18481 9276
rect 18537 9274 18561 9276
rect 18617 9274 18623 9276
rect 18377 9222 18379 9274
rect 18559 9222 18561 9274
rect 18315 9220 18321 9222
rect 18377 9220 18401 9222
rect 18457 9220 18481 9222
rect 18537 9220 18561 9222
rect 18617 9220 18623 9222
rect 18315 9211 18623 9220
rect 25261 9276 25569 9285
rect 25261 9274 25267 9276
rect 25323 9274 25347 9276
rect 25403 9274 25427 9276
rect 25483 9274 25507 9276
rect 25563 9274 25569 9276
rect 25323 9222 25325 9274
rect 25505 9222 25507 9274
rect 25261 9220 25267 9222
rect 25323 9220 25347 9222
rect 25403 9220 25427 9222
rect 25483 9220 25507 9222
rect 25563 9220 25569 9222
rect 25261 9211 25569 9220
rect 28356 9104 28408 9110
rect 28354 9072 28356 9081
rect 28408 9072 28410 9081
rect 28354 9007 28410 9016
rect 21788 8732 22096 8741
rect 21788 8730 21794 8732
rect 21850 8730 21874 8732
rect 21930 8730 21954 8732
rect 22010 8730 22034 8732
rect 22090 8730 22096 8732
rect 21850 8678 21852 8730
rect 22032 8678 22034 8730
rect 21788 8676 21794 8678
rect 21850 8676 21874 8678
rect 21930 8676 21954 8678
rect 22010 8676 22034 8678
rect 22090 8676 22096 8678
rect 21788 8667 22096 8676
rect 28734 8732 29042 8741
rect 28734 8730 28740 8732
rect 28796 8730 28820 8732
rect 28876 8730 28900 8732
rect 28956 8730 28980 8732
rect 29036 8730 29042 8732
rect 28796 8678 28798 8730
rect 28978 8678 28980 8730
rect 28734 8676 28740 8678
rect 28796 8676 28820 8678
rect 28876 8676 28900 8678
rect 28956 8676 28980 8678
rect 29036 8676 29042 8678
rect 28734 8667 29042 8676
rect 18315 8188 18623 8197
rect 18315 8186 18321 8188
rect 18377 8186 18401 8188
rect 18457 8186 18481 8188
rect 18537 8186 18561 8188
rect 18617 8186 18623 8188
rect 18377 8134 18379 8186
rect 18559 8134 18561 8186
rect 18315 8132 18321 8134
rect 18377 8132 18401 8134
rect 18457 8132 18481 8134
rect 18537 8132 18561 8134
rect 18617 8132 18623 8134
rect 18315 8123 18623 8132
rect 25261 8188 25569 8197
rect 25261 8186 25267 8188
rect 25323 8186 25347 8188
rect 25403 8186 25427 8188
rect 25483 8186 25507 8188
rect 25563 8186 25569 8188
rect 25323 8134 25325 8186
rect 25505 8134 25507 8186
rect 25261 8132 25267 8134
rect 25323 8132 25347 8134
rect 25403 8132 25427 8134
rect 25483 8132 25507 8134
rect 25563 8132 25569 8134
rect 25261 8123 25569 8132
rect 28356 7880 28408 7886
rect 28356 7822 28408 7828
rect 21788 7644 22096 7653
rect 21788 7642 21794 7644
rect 21850 7642 21874 7644
rect 21930 7642 21954 7644
rect 22010 7642 22034 7644
rect 22090 7642 22096 7644
rect 21850 7590 21852 7642
rect 22032 7590 22034 7642
rect 21788 7588 21794 7590
rect 21850 7588 21874 7590
rect 21930 7588 21954 7590
rect 22010 7588 22034 7590
rect 22090 7588 22096 7590
rect 21788 7579 22096 7588
rect 28368 7449 28396 7822
rect 28734 7644 29042 7653
rect 28734 7642 28740 7644
rect 28796 7642 28820 7644
rect 28876 7642 28900 7644
rect 28956 7642 28980 7644
rect 29036 7642 29042 7644
rect 28796 7590 28798 7642
rect 28978 7590 28980 7642
rect 28734 7588 28740 7590
rect 28796 7588 28820 7590
rect 28876 7588 28900 7590
rect 28956 7588 28980 7590
rect 29036 7588 29042 7590
rect 28734 7579 29042 7588
rect 28354 7440 28410 7449
rect 28354 7375 28410 7384
rect 18315 7100 18623 7109
rect 18315 7098 18321 7100
rect 18377 7098 18401 7100
rect 18457 7098 18481 7100
rect 18537 7098 18561 7100
rect 18617 7098 18623 7100
rect 18377 7046 18379 7098
rect 18559 7046 18561 7098
rect 18315 7044 18321 7046
rect 18377 7044 18401 7046
rect 18457 7044 18481 7046
rect 18537 7044 18561 7046
rect 18617 7044 18623 7046
rect 18315 7035 18623 7044
rect 25261 7100 25569 7109
rect 25261 7098 25267 7100
rect 25323 7098 25347 7100
rect 25403 7098 25427 7100
rect 25483 7098 25507 7100
rect 25563 7098 25569 7100
rect 25323 7046 25325 7098
rect 25505 7046 25507 7098
rect 25261 7044 25267 7046
rect 25323 7044 25347 7046
rect 25403 7044 25427 7046
rect 25483 7044 25507 7046
rect 25563 7044 25569 7046
rect 25261 7035 25569 7044
rect 28356 6792 28408 6798
rect 28354 6760 28356 6769
rect 28408 6760 28410 6769
rect 28354 6695 28410 6704
rect 21788 6556 22096 6565
rect 21788 6554 21794 6556
rect 21850 6554 21874 6556
rect 21930 6554 21954 6556
rect 22010 6554 22034 6556
rect 22090 6554 22096 6556
rect 21850 6502 21852 6554
rect 22032 6502 22034 6554
rect 21788 6500 21794 6502
rect 21850 6500 21874 6502
rect 21930 6500 21954 6502
rect 22010 6500 22034 6502
rect 22090 6500 22096 6502
rect 21788 6491 22096 6500
rect 28734 6556 29042 6565
rect 28734 6554 28740 6556
rect 28796 6554 28820 6556
rect 28876 6554 28900 6556
rect 28956 6554 28980 6556
rect 29036 6554 29042 6556
rect 28796 6502 28798 6554
rect 28978 6502 28980 6554
rect 28734 6500 28740 6502
rect 28796 6500 28820 6502
rect 28876 6500 28900 6502
rect 28956 6500 28980 6502
rect 29036 6500 29042 6502
rect 28734 6491 29042 6500
rect 18315 6012 18623 6021
rect 18315 6010 18321 6012
rect 18377 6010 18401 6012
rect 18457 6010 18481 6012
rect 18537 6010 18561 6012
rect 18617 6010 18623 6012
rect 18377 5958 18379 6010
rect 18559 5958 18561 6010
rect 18315 5956 18321 5958
rect 18377 5956 18401 5958
rect 18457 5956 18481 5958
rect 18537 5956 18561 5958
rect 18617 5956 18623 5958
rect 18315 5947 18623 5956
rect 25261 6012 25569 6021
rect 25261 6010 25267 6012
rect 25323 6010 25347 6012
rect 25403 6010 25427 6012
rect 25483 6010 25507 6012
rect 25563 6010 25569 6012
rect 25323 5958 25325 6010
rect 25505 5958 25507 6010
rect 25261 5956 25267 5958
rect 25323 5956 25347 5958
rect 25403 5956 25427 5958
rect 25483 5956 25507 5958
rect 25563 5956 25569 5958
rect 25261 5947 25569 5956
rect 28356 5704 28408 5710
rect 28354 5672 28356 5681
rect 28408 5672 28410 5681
rect 28354 5607 28410 5616
rect 21788 5468 22096 5477
rect 21788 5466 21794 5468
rect 21850 5466 21874 5468
rect 21930 5466 21954 5468
rect 22010 5466 22034 5468
rect 22090 5466 22096 5468
rect 21850 5414 21852 5466
rect 22032 5414 22034 5466
rect 21788 5412 21794 5414
rect 21850 5412 21874 5414
rect 21930 5412 21954 5414
rect 22010 5412 22034 5414
rect 22090 5412 22096 5414
rect 21788 5403 22096 5412
rect 28734 5468 29042 5477
rect 28734 5466 28740 5468
rect 28796 5466 28820 5468
rect 28876 5466 28900 5468
rect 28956 5466 28980 5468
rect 29036 5466 29042 5468
rect 28796 5414 28798 5466
rect 28978 5414 28980 5466
rect 28734 5412 28740 5414
rect 28796 5412 28820 5414
rect 28876 5412 28900 5414
rect 28956 5412 28980 5414
rect 29036 5412 29042 5414
rect 28734 5403 29042 5412
rect 28356 5024 28408 5030
rect 28356 4966 28408 4972
rect 18315 4924 18623 4933
rect 18315 4922 18321 4924
rect 18377 4922 18401 4924
rect 18457 4922 18481 4924
rect 18537 4922 18561 4924
rect 18617 4922 18623 4924
rect 18377 4870 18379 4922
rect 18559 4870 18561 4922
rect 18315 4868 18321 4870
rect 18377 4868 18401 4870
rect 18457 4868 18481 4870
rect 18537 4868 18561 4870
rect 18617 4868 18623 4870
rect 18315 4859 18623 4868
rect 25261 4924 25569 4933
rect 25261 4922 25267 4924
rect 25323 4922 25347 4924
rect 25403 4922 25427 4924
rect 25483 4922 25507 4924
rect 25563 4922 25569 4924
rect 25323 4870 25325 4922
rect 25505 4870 25507 4922
rect 25261 4868 25267 4870
rect 25323 4868 25347 4870
rect 25403 4868 25427 4870
rect 25483 4868 25507 4870
rect 25563 4868 25569 4870
rect 25261 4859 25569 4868
rect 28368 4729 28396 4966
rect 28354 4720 28410 4729
rect 28354 4655 28410 4664
rect 28356 4480 28408 4486
rect 28356 4422 28408 4428
rect 21788 4380 22096 4389
rect 21788 4378 21794 4380
rect 21850 4378 21874 4380
rect 21930 4378 21954 4380
rect 22010 4378 22034 4380
rect 22090 4378 22096 4380
rect 21850 4326 21852 4378
rect 22032 4326 22034 4378
rect 21788 4324 21794 4326
rect 21850 4324 21874 4326
rect 21930 4324 21954 4326
rect 22010 4324 22034 4326
rect 22090 4324 22096 4326
rect 21788 4315 22096 4324
rect 28368 4078 28396 4422
rect 28734 4380 29042 4389
rect 28734 4378 28740 4380
rect 28796 4378 28820 4380
rect 28876 4378 28900 4380
rect 28956 4378 28980 4380
rect 29036 4378 29042 4380
rect 28796 4326 28798 4378
rect 28978 4326 28980 4378
rect 28734 4324 28740 4326
rect 28796 4324 28820 4326
rect 28876 4324 28900 4326
rect 28956 4324 28980 4326
rect 29036 4324 29042 4326
rect 28734 4315 29042 4324
rect 17132 4072 17184 4078
rect 28356 4072 28408 4078
rect 17132 4014 17184 4020
rect 28354 4040 28356 4049
rect 28408 4040 28410 4049
rect 28354 3975 28410 3984
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 1596 3777 1624 3878
rect 4423 3836 4731 3845
rect 4423 3834 4429 3836
rect 4485 3834 4509 3836
rect 4565 3834 4589 3836
rect 4645 3834 4669 3836
rect 4725 3834 4731 3836
rect 4485 3782 4487 3834
rect 4667 3782 4669 3834
rect 4423 3780 4429 3782
rect 4485 3780 4509 3782
rect 4565 3780 4589 3782
rect 4645 3780 4669 3782
rect 4725 3780 4731 3782
rect 1582 3768 1638 3777
rect 4423 3771 4731 3780
rect 11369 3836 11677 3845
rect 11369 3834 11375 3836
rect 11431 3834 11455 3836
rect 11511 3834 11535 3836
rect 11591 3834 11615 3836
rect 11671 3834 11677 3836
rect 11431 3782 11433 3834
rect 11613 3782 11615 3834
rect 11369 3780 11375 3782
rect 11431 3780 11455 3782
rect 11511 3780 11535 3782
rect 11591 3780 11615 3782
rect 11671 3780 11677 3782
rect 11369 3771 11677 3780
rect 18315 3836 18623 3845
rect 18315 3834 18321 3836
rect 18377 3834 18401 3836
rect 18457 3834 18481 3836
rect 18537 3834 18561 3836
rect 18617 3834 18623 3836
rect 18377 3782 18379 3834
rect 18559 3782 18561 3834
rect 18315 3780 18321 3782
rect 18377 3780 18401 3782
rect 18457 3780 18481 3782
rect 18537 3780 18561 3782
rect 18617 3780 18623 3782
rect 18315 3771 18623 3780
rect 25261 3836 25569 3845
rect 25261 3834 25267 3836
rect 25323 3834 25347 3836
rect 25403 3834 25427 3836
rect 25483 3834 25507 3836
rect 25563 3834 25569 3836
rect 25323 3782 25325 3834
rect 25505 3782 25507 3834
rect 25261 3780 25267 3782
rect 25323 3780 25347 3782
rect 25403 3780 25427 3782
rect 25483 3780 25507 3782
rect 25563 3780 25569 3782
rect 25261 3771 25569 3780
rect 1582 3703 1638 3712
rect 28356 3664 28408 3670
rect 28354 3632 28356 3641
rect 28408 3632 28410 3641
rect 28354 3567 28410 3576
rect 1584 3528 1636 3534
rect 1584 3470 1636 3476
rect 1596 3097 1624 3470
rect 7896 3292 8204 3301
rect 7896 3290 7902 3292
rect 7958 3290 7982 3292
rect 8038 3290 8062 3292
rect 8118 3290 8142 3292
rect 8198 3290 8204 3292
rect 7958 3238 7960 3290
rect 8140 3238 8142 3290
rect 7896 3236 7902 3238
rect 7958 3236 7982 3238
rect 8038 3236 8062 3238
rect 8118 3236 8142 3238
rect 8198 3236 8204 3238
rect 7896 3227 8204 3236
rect 14842 3292 15150 3301
rect 14842 3290 14848 3292
rect 14904 3290 14928 3292
rect 14984 3290 15008 3292
rect 15064 3290 15088 3292
rect 15144 3290 15150 3292
rect 14904 3238 14906 3290
rect 15086 3238 15088 3290
rect 14842 3236 14848 3238
rect 14904 3236 14928 3238
rect 14984 3236 15008 3238
rect 15064 3236 15088 3238
rect 15144 3236 15150 3238
rect 14842 3227 15150 3236
rect 21788 3292 22096 3301
rect 21788 3290 21794 3292
rect 21850 3290 21874 3292
rect 21930 3290 21954 3292
rect 22010 3290 22034 3292
rect 22090 3290 22096 3292
rect 21850 3238 21852 3290
rect 22032 3238 22034 3290
rect 21788 3236 21794 3238
rect 21850 3236 21874 3238
rect 21930 3236 21954 3238
rect 22010 3236 22034 3238
rect 22090 3236 22096 3238
rect 21788 3227 22096 3236
rect 28734 3292 29042 3301
rect 28734 3290 28740 3292
rect 28796 3290 28820 3292
rect 28876 3290 28900 3292
rect 28956 3290 28980 3292
rect 29036 3290 29042 3292
rect 28796 3238 28798 3290
rect 28978 3238 28980 3290
rect 28734 3236 28740 3238
rect 28796 3236 28820 3238
rect 28876 3236 28900 3238
rect 28956 3236 28980 3238
rect 29036 3236 29042 3238
rect 28734 3227 29042 3236
rect 1582 3088 1638 3097
rect 1582 3023 1638 3032
rect 28356 2848 28408 2854
rect 28356 2790 28408 2796
rect 4423 2748 4731 2757
rect 4423 2746 4429 2748
rect 4485 2746 4509 2748
rect 4565 2746 4589 2748
rect 4645 2746 4669 2748
rect 4725 2746 4731 2748
rect 4485 2694 4487 2746
rect 4667 2694 4669 2746
rect 4423 2692 4429 2694
rect 4485 2692 4509 2694
rect 4565 2692 4589 2694
rect 4645 2692 4669 2694
rect 4725 2692 4731 2694
rect 4423 2683 4731 2692
rect 11369 2748 11677 2757
rect 11369 2746 11375 2748
rect 11431 2746 11455 2748
rect 11511 2746 11535 2748
rect 11591 2746 11615 2748
rect 11671 2746 11677 2748
rect 11431 2694 11433 2746
rect 11613 2694 11615 2746
rect 11369 2692 11375 2694
rect 11431 2692 11455 2694
rect 11511 2692 11535 2694
rect 11591 2692 11615 2694
rect 11671 2692 11677 2694
rect 11369 2683 11677 2692
rect 18315 2748 18623 2757
rect 18315 2746 18321 2748
rect 18377 2746 18401 2748
rect 18457 2746 18481 2748
rect 18537 2746 18561 2748
rect 18617 2746 18623 2748
rect 18377 2694 18379 2746
rect 18559 2694 18561 2746
rect 18315 2692 18321 2694
rect 18377 2692 18401 2694
rect 18457 2692 18481 2694
rect 18537 2692 18561 2694
rect 18617 2692 18623 2694
rect 18315 2683 18623 2692
rect 25261 2748 25569 2757
rect 25261 2746 25267 2748
rect 25323 2746 25347 2748
rect 25403 2746 25427 2748
rect 25483 2746 25507 2748
rect 25563 2746 25569 2748
rect 25323 2694 25325 2746
rect 25505 2694 25507 2746
rect 25261 2692 25267 2694
rect 25323 2692 25347 2694
rect 25403 2692 25427 2694
rect 25483 2692 25507 2694
rect 25563 2692 25569 2694
rect 25261 2683 25569 2692
rect 28368 2689 28396 2790
rect 28354 2680 28410 2689
rect 28354 2615 28410 2624
rect 7896 2204 8204 2213
rect 7896 2202 7902 2204
rect 7958 2202 7982 2204
rect 8038 2202 8062 2204
rect 8118 2202 8142 2204
rect 8198 2202 8204 2204
rect 7958 2150 7960 2202
rect 8140 2150 8142 2202
rect 7896 2148 7902 2150
rect 7958 2148 7982 2150
rect 8038 2148 8062 2150
rect 8118 2148 8142 2150
rect 8198 2148 8204 2150
rect 7896 2139 8204 2148
rect 14842 2204 15150 2213
rect 14842 2202 14848 2204
rect 14904 2202 14928 2204
rect 14984 2202 15008 2204
rect 15064 2202 15088 2204
rect 15144 2202 15150 2204
rect 14904 2150 14906 2202
rect 15086 2150 15088 2202
rect 14842 2148 14848 2150
rect 14904 2148 14928 2150
rect 14984 2148 15008 2150
rect 15064 2148 15088 2150
rect 15144 2148 15150 2150
rect 14842 2139 15150 2148
rect 21788 2204 22096 2213
rect 21788 2202 21794 2204
rect 21850 2202 21874 2204
rect 21930 2202 21954 2204
rect 22010 2202 22034 2204
rect 22090 2202 22096 2204
rect 21850 2150 21852 2202
rect 22032 2150 22034 2202
rect 21788 2148 21794 2150
rect 21850 2148 21874 2150
rect 21930 2148 21954 2150
rect 22010 2148 22034 2150
rect 22090 2148 22096 2150
rect 21788 2139 22096 2148
rect 28734 2204 29042 2213
rect 28734 2202 28740 2204
rect 28796 2202 28820 2204
rect 28876 2202 28900 2204
rect 28956 2202 28980 2204
rect 29036 2202 29042 2204
rect 28796 2150 28798 2202
rect 28978 2150 28980 2202
rect 28734 2148 28740 2150
rect 28796 2148 28820 2150
rect 28876 2148 28900 2150
rect 28956 2148 28980 2150
rect 29036 2148 29042 2150
rect 28734 2139 29042 2148
<< via2 >>
rect 1674 28192 1730 28248
rect 1582 26152 1638 26208
rect 2870 30232 2926 30288
rect 2318 30096 2374 30152
rect 2594 29572 2650 29608
rect 2594 29552 2596 29572
rect 2596 29552 2648 29572
rect 2648 29552 2650 29572
rect 2042 27920 2098 27976
rect 2226 27376 2282 27432
rect 2778 27512 2834 27568
rect 2594 26288 2650 26344
rect 2318 26188 2320 26208
rect 2320 26188 2372 26208
rect 2372 26188 2374 26208
rect 2318 26152 2374 26188
rect 2318 25472 2374 25528
rect 2962 29416 3018 29472
rect 3238 28600 3294 28656
rect 3238 26968 3294 27024
rect 3238 25744 3294 25800
rect 3698 26832 3754 26888
rect 3790 26016 3846 26072
rect 4429 31034 4485 31036
rect 4509 31034 4565 31036
rect 4589 31034 4645 31036
rect 4669 31034 4725 31036
rect 4429 30982 4475 31034
rect 4475 30982 4485 31034
rect 4509 30982 4539 31034
rect 4539 30982 4551 31034
rect 4551 30982 4565 31034
rect 4589 30982 4603 31034
rect 4603 30982 4615 31034
rect 4615 30982 4645 31034
rect 4669 30982 4679 31034
rect 4679 30982 4725 31034
rect 4429 30980 4485 30982
rect 4509 30980 4565 30982
rect 4589 30980 4645 30982
rect 4669 30980 4725 30982
rect 3974 28600 4030 28656
rect 4158 28600 4214 28656
rect 3330 24792 3386 24848
rect 4429 29946 4485 29948
rect 4509 29946 4565 29948
rect 4589 29946 4645 29948
rect 4669 29946 4725 29948
rect 4429 29894 4475 29946
rect 4475 29894 4485 29946
rect 4509 29894 4539 29946
rect 4539 29894 4551 29946
rect 4551 29894 4565 29946
rect 4589 29894 4603 29946
rect 4603 29894 4615 29946
rect 4615 29894 4645 29946
rect 4669 29894 4679 29946
rect 4679 29894 4725 29946
rect 4429 29892 4485 29894
rect 4509 29892 4565 29894
rect 4589 29892 4645 29894
rect 4669 29892 4725 29894
rect 4429 28858 4485 28860
rect 4509 28858 4565 28860
rect 4589 28858 4645 28860
rect 4669 28858 4725 28860
rect 4429 28806 4475 28858
rect 4475 28806 4485 28858
rect 4509 28806 4539 28858
rect 4539 28806 4551 28858
rect 4551 28806 4565 28858
rect 4589 28806 4603 28858
rect 4603 28806 4615 28858
rect 4615 28806 4645 28858
rect 4669 28806 4679 28858
rect 4679 28806 4725 28858
rect 4429 28804 4485 28806
rect 4509 28804 4565 28806
rect 4589 28804 4645 28806
rect 4669 28804 4725 28806
rect 4429 27770 4485 27772
rect 4509 27770 4565 27772
rect 4589 27770 4645 27772
rect 4669 27770 4725 27772
rect 4429 27718 4475 27770
rect 4475 27718 4485 27770
rect 4509 27718 4539 27770
rect 4539 27718 4551 27770
rect 4551 27718 4565 27770
rect 4589 27718 4603 27770
rect 4603 27718 4615 27770
rect 4615 27718 4645 27770
rect 4669 27718 4679 27770
rect 4679 27718 4725 27770
rect 4429 27716 4485 27718
rect 4509 27716 4565 27718
rect 4589 27716 4645 27718
rect 4669 27716 4725 27718
rect 4710 27104 4766 27160
rect 4429 26682 4485 26684
rect 4509 26682 4565 26684
rect 4589 26682 4645 26684
rect 4669 26682 4725 26684
rect 4429 26630 4475 26682
rect 4475 26630 4485 26682
rect 4509 26630 4539 26682
rect 4539 26630 4551 26682
rect 4551 26630 4565 26682
rect 4589 26630 4603 26682
rect 4603 26630 4615 26682
rect 4615 26630 4645 26682
rect 4669 26630 4679 26682
rect 4679 26630 4725 26682
rect 4429 26628 4485 26630
rect 4509 26628 4565 26630
rect 4589 26628 4645 26630
rect 4669 26628 4725 26630
rect 4434 26460 4436 26480
rect 4436 26460 4488 26480
rect 4488 26460 4490 26480
rect 4434 26424 4490 26460
rect 4429 25594 4485 25596
rect 4509 25594 4565 25596
rect 4589 25594 4645 25596
rect 4669 25594 4725 25596
rect 4429 25542 4475 25594
rect 4475 25542 4485 25594
rect 4509 25542 4539 25594
rect 4539 25542 4551 25594
rect 4551 25542 4565 25594
rect 4589 25542 4603 25594
rect 4603 25542 4615 25594
rect 4615 25542 4645 25594
rect 4669 25542 4679 25594
rect 4679 25542 4725 25594
rect 4429 25540 4485 25542
rect 4509 25540 4565 25542
rect 4589 25540 4645 25542
rect 4669 25540 4725 25542
rect 4250 25200 4306 25256
rect 4429 24506 4485 24508
rect 4509 24506 4565 24508
rect 4589 24506 4645 24508
rect 4669 24506 4725 24508
rect 4429 24454 4475 24506
rect 4475 24454 4485 24506
rect 4509 24454 4539 24506
rect 4539 24454 4551 24506
rect 4551 24454 4565 24506
rect 4589 24454 4603 24506
rect 4603 24454 4615 24506
rect 4615 24454 4645 24506
rect 4669 24454 4679 24506
rect 4679 24454 4725 24506
rect 4429 24452 4485 24454
rect 4509 24452 4565 24454
rect 4589 24452 4645 24454
rect 4669 24452 4725 24454
rect 5446 31340 5502 31376
rect 5446 31320 5448 31340
rect 5448 31320 5500 31340
rect 5500 31320 5502 31340
rect 6090 30268 6092 30288
rect 6092 30268 6144 30288
rect 6144 30268 6146 30288
rect 6090 30232 6146 30268
rect 5262 25880 5318 25936
rect 5722 26696 5778 26752
rect 5538 26288 5594 26344
rect 5998 29144 6054 29200
rect 6642 31184 6698 31240
rect 6734 30368 6790 30424
rect 6274 27104 6330 27160
rect 5998 26152 6054 26208
rect 6458 27396 6514 27432
rect 6458 27376 6460 27396
rect 6460 27376 6512 27396
rect 6512 27376 6514 27396
rect 6366 26696 6422 26752
rect 5170 24928 5226 24984
rect 1582 24148 1584 24168
rect 1584 24148 1636 24168
rect 1636 24148 1638 24168
rect 1582 24112 1638 24148
rect 6642 26560 6698 26616
rect 6458 25472 6514 25528
rect 7010 30268 7012 30288
rect 7012 30268 7064 30288
rect 7064 30268 7066 30288
rect 7010 30232 7066 30268
rect 7902 31578 7958 31580
rect 7982 31578 8038 31580
rect 8062 31578 8118 31580
rect 8142 31578 8198 31580
rect 7902 31526 7948 31578
rect 7948 31526 7958 31578
rect 7982 31526 8012 31578
rect 8012 31526 8024 31578
rect 8024 31526 8038 31578
rect 8062 31526 8076 31578
rect 8076 31526 8088 31578
rect 8088 31526 8118 31578
rect 8142 31526 8152 31578
rect 8152 31526 8198 31578
rect 7902 31524 7958 31526
rect 7982 31524 8038 31526
rect 8062 31524 8118 31526
rect 8142 31524 8198 31526
rect 7562 30776 7618 30832
rect 7194 30640 7250 30696
rect 7102 28872 7158 28928
rect 7194 26016 7250 26072
rect 7902 30490 7958 30492
rect 7982 30490 8038 30492
rect 8062 30490 8118 30492
rect 8142 30490 8198 30492
rect 7902 30438 7948 30490
rect 7948 30438 7958 30490
rect 7982 30438 8012 30490
rect 8012 30438 8024 30490
rect 8024 30438 8038 30490
rect 8062 30438 8076 30490
rect 8076 30438 8088 30490
rect 8088 30438 8118 30490
rect 8142 30438 8152 30490
rect 8152 30438 8198 30490
rect 7902 30436 7958 30438
rect 7982 30436 8038 30438
rect 8062 30436 8118 30438
rect 8142 30436 8198 30438
rect 7902 29402 7958 29404
rect 7982 29402 8038 29404
rect 8062 29402 8118 29404
rect 8142 29402 8198 29404
rect 7902 29350 7948 29402
rect 7948 29350 7958 29402
rect 7982 29350 8012 29402
rect 8012 29350 8024 29402
rect 8024 29350 8038 29402
rect 8062 29350 8076 29402
rect 8076 29350 8088 29402
rect 8088 29350 8118 29402
rect 8142 29350 8152 29402
rect 8152 29350 8198 29402
rect 7902 29348 7958 29350
rect 7982 29348 8038 29350
rect 8062 29348 8118 29350
rect 8142 29348 8198 29350
rect 7562 29044 7564 29064
rect 7564 29044 7616 29064
rect 7616 29044 7618 29064
rect 7562 29008 7618 29044
rect 8390 29028 8446 29064
rect 8390 29008 8392 29028
rect 8392 29008 8444 29028
rect 8444 29008 8446 29028
rect 7654 26560 7710 26616
rect 7562 25472 7618 25528
rect 7470 25336 7526 25392
rect 7562 24928 7618 24984
rect 7902 28314 7958 28316
rect 7982 28314 8038 28316
rect 8062 28314 8118 28316
rect 8142 28314 8198 28316
rect 7902 28262 7948 28314
rect 7948 28262 7958 28314
rect 7982 28262 8012 28314
rect 8012 28262 8024 28314
rect 8024 28262 8038 28314
rect 8062 28262 8076 28314
rect 8076 28262 8088 28314
rect 8088 28262 8118 28314
rect 8142 28262 8152 28314
rect 8152 28262 8198 28314
rect 7902 28260 7958 28262
rect 7982 28260 8038 28262
rect 8062 28260 8118 28262
rect 8142 28260 8198 28262
rect 7902 27226 7958 27228
rect 7982 27226 8038 27228
rect 8062 27226 8118 27228
rect 8142 27226 8198 27228
rect 7902 27174 7948 27226
rect 7948 27174 7958 27226
rect 7982 27174 8012 27226
rect 8012 27174 8024 27226
rect 8024 27174 8038 27226
rect 8062 27174 8076 27226
rect 8076 27174 8088 27226
rect 8088 27174 8118 27226
rect 8142 27174 8152 27226
rect 8152 27174 8198 27226
rect 7902 27172 7958 27174
rect 7982 27172 8038 27174
rect 8062 27172 8118 27174
rect 8142 27172 8198 27174
rect 7902 26138 7958 26140
rect 7982 26138 8038 26140
rect 8062 26138 8118 26140
rect 8142 26138 8198 26140
rect 7902 26086 7948 26138
rect 7948 26086 7958 26138
rect 7982 26086 8012 26138
rect 8012 26086 8024 26138
rect 8024 26086 8038 26138
rect 8062 26086 8076 26138
rect 8076 26086 8088 26138
rect 8088 26086 8118 26138
rect 8142 26086 8152 26138
rect 8152 26086 8198 26138
rect 7902 26084 7958 26086
rect 7982 26084 8038 26086
rect 8062 26084 8118 26086
rect 8142 26084 8198 26086
rect 7838 25336 7894 25392
rect 7902 25050 7958 25052
rect 7982 25050 8038 25052
rect 8062 25050 8118 25052
rect 8142 25050 8198 25052
rect 7902 24998 7948 25050
rect 7948 24998 7958 25050
rect 7982 24998 8012 25050
rect 8012 24998 8024 25050
rect 8024 24998 8038 25050
rect 8062 24998 8076 25050
rect 8076 24998 8088 25050
rect 8088 24998 8118 25050
rect 8142 24998 8152 25050
rect 8152 24998 8198 25050
rect 7902 24996 7958 24998
rect 7982 24996 8038 24998
rect 8062 24996 8118 24998
rect 8142 24996 8198 24998
rect 8666 28600 8722 28656
rect 8758 27376 8814 27432
rect 8390 26460 8392 26480
rect 8392 26460 8444 26480
rect 8444 26460 8446 26480
rect 8390 26424 8446 26460
rect 8758 26560 8814 26616
rect 8942 29008 8998 29064
rect 9034 26968 9090 27024
rect 7902 23962 7958 23964
rect 7982 23962 8038 23964
rect 8062 23962 8118 23964
rect 8142 23962 8198 23964
rect 7902 23910 7948 23962
rect 7948 23910 7958 23962
rect 7982 23910 8012 23962
rect 8012 23910 8024 23962
rect 8024 23910 8038 23962
rect 8062 23910 8076 23962
rect 8076 23910 8088 23962
rect 8088 23910 8118 23962
rect 8142 23910 8152 23962
rect 8152 23910 8198 23962
rect 7902 23908 7958 23910
rect 7982 23908 8038 23910
rect 8062 23908 8118 23910
rect 8142 23908 8198 23910
rect 11794 31048 11850 31104
rect 11375 31034 11431 31036
rect 11455 31034 11511 31036
rect 11535 31034 11591 31036
rect 11615 31034 11671 31036
rect 11375 30982 11421 31034
rect 11421 30982 11431 31034
rect 11455 30982 11485 31034
rect 11485 30982 11497 31034
rect 11497 30982 11511 31034
rect 11535 30982 11549 31034
rect 11549 30982 11561 31034
rect 11561 30982 11591 31034
rect 11615 30982 11625 31034
rect 11625 30982 11671 31034
rect 11375 30980 11431 30982
rect 11455 30980 11511 30982
rect 11535 30980 11591 30982
rect 11615 30980 11671 30982
rect 9678 30232 9734 30288
rect 8666 24656 8722 24712
rect 10230 29280 10286 29336
rect 9862 28872 9918 28928
rect 9678 28056 9734 28112
rect 9954 28192 10010 28248
rect 9862 26016 9918 26072
rect 9770 25356 9826 25392
rect 9770 25336 9772 25356
rect 9772 25336 9824 25356
rect 9824 25336 9826 25356
rect 10322 26152 10378 26208
rect 10414 26016 10470 26072
rect 11150 30504 11206 30560
rect 9586 24692 9588 24712
rect 9588 24692 9640 24712
rect 9640 24692 9642 24712
rect 9586 24656 9642 24692
rect 1582 23468 1584 23488
rect 1584 23468 1636 23488
rect 1636 23468 1638 23488
rect 1582 23432 1638 23468
rect 4429 23418 4485 23420
rect 4509 23418 4565 23420
rect 4589 23418 4645 23420
rect 4669 23418 4725 23420
rect 4429 23366 4475 23418
rect 4475 23366 4485 23418
rect 4509 23366 4539 23418
rect 4539 23366 4551 23418
rect 4551 23366 4565 23418
rect 4589 23366 4603 23418
rect 4603 23366 4615 23418
rect 4615 23366 4645 23418
rect 4669 23366 4679 23418
rect 4679 23366 4725 23418
rect 4429 23364 4485 23366
rect 4509 23364 4565 23366
rect 4589 23364 4645 23366
rect 4669 23364 4725 23366
rect 10598 25200 10654 25256
rect 10966 27512 11022 27568
rect 11150 29144 11206 29200
rect 11794 30640 11850 30696
rect 11794 30232 11850 30288
rect 11375 29946 11431 29948
rect 11455 29946 11511 29948
rect 11535 29946 11591 29948
rect 11615 29946 11671 29948
rect 11375 29894 11421 29946
rect 11421 29894 11431 29946
rect 11455 29894 11485 29946
rect 11485 29894 11497 29946
rect 11497 29894 11511 29946
rect 11535 29894 11549 29946
rect 11549 29894 11561 29946
rect 11561 29894 11591 29946
rect 11615 29894 11625 29946
rect 11625 29894 11671 29946
rect 11375 29892 11431 29894
rect 11455 29892 11511 29894
rect 11535 29892 11591 29894
rect 11615 29892 11671 29894
rect 11375 28858 11431 28860
rect 11455 28858 11511 28860
rect 11535 28858 11591 28860
rect 11615 28858 11671 28860
rect 11375 28806 11421 28858
rect 11421 28806 11431 28858
rect 11455 28806 11485 28858
rect 11485 28806 11497 28858
rect 11497 28806 11511 28858
rect 11535 28806 11549 28858
rect 11549 28806 11561 28858
rect 11561 28806 11591 28858
rect 11615 28806 11625 28858
rect 11625 28806 11671 28858
rect 11375 28804 11431 28806
rect 11455 28804 11511 28806
rect 11535 28804 11591 28806
rect 11615 28804 11671 28806
rect 12162 30640 12218 30696
rect 12438 29960 12494 30016
rect 12070 29688 12126 29744
rect 11794 28736 11850 28792
rect 11794 28600 11850 28656
rect 11375 27770 11431 27772
rect 11455 27770 11511 27772
rect 11535 27770 11591 27772
rect 11615 27770 11671 27772
rect 11375 27718 11421 27770
rect 11421 27718 11431 27770
rect 11455 27718 11485 27770
rect 11485 27718 11497 27770
rect 11497 27718 11511 27770
rect 11535 27718 11549 27770
rect 11549 27718 11561 27770
rect 11561 27718 11591 27770
rect 11615 27718 11625 27770
rect 11625 27718 11671 27770
rect 11375 27716 11431 27718
rect 11455 27716 11511 27718
rect 11535 27716 11591 27718
rect 11615 27716 11671 27718
rect 11375 26682 11431 26684
rect 11455 26682 11511 26684
rect 11535 26682 11591 26684
rect 11615 26682 11671 26684
rect 11375 26630 11421 26682
rect 11421 26630 11431 26682
rect 11455 26630 11485 26682
rect 11485 26630 11497 26682
rect 11497 26630 11511 26682
rect 11535 26630 11549 26682
rect 11549 26630 11561 26682
rect 11561 26630 11591 26682
rect 11615 26630 11625 26682
rect 11625 26630 11671 26682
rect 11375 26628 11431 26630
rect 11455 26628 11511 26630
rect 11535 26628 11591 26630
rect 11615 26628 11671 26630
rect 11702 25916 11704 25936
rect 11704 25916 11756 25936
rect 11756 25916 11758 25936
rect 11702 25880 11758 25916
rect 11375 25594 11431 25596
rect 11455 25594 11511 25596
rect 11535 25594 11591 25596
rect 11615 25594 11671 25596
rect 11375 25542 11421 25594
rect 11421 25542 11431 25594
rect 11455 25542 11485 25594
rect 11485 25542 11497 25594
rect 11497 25542 11511 25594
rect 11535 25542 11549 25594
rect 11549 25542 11561 25594
rect 11561 25542 11591 25594
rect 11615 25542 11625 25594
rect 11625 25542 11671 25594
rect 11375 25540 11431 25542
rect 11455 25540 11511 25542
rect 11535 25540 11591 25542
rect 11615 25540 11671 25542
rect 11058 25336 11114 25392
rect 11702 24792 11758 24848
rect 11375 24506 11431 24508
rect 11455 24506 11511 24508
rect 11535 24506 11591 24508
rect 11615 24506 11671 24508
rect 11375 24454 11421 24506
rect 11421 24454 11431 24506
rect 11455 24454 11485 24506
rect 11485 24454 11497 24506
rect 11497 24454 11511 24506
rect 11535 24454 11549 24506
rect 11549 24454 11561 24506
rect 11561 24454 11591 24506
rect 11615 24454 11625 24506
rect 11625 24454 11671 24506
rect 11375 24452 11431 24454
rect 11455 24452 11511 24454
rect 11535 24452 11591 24454
rect 11615 24452 11671 24454
rect 12254 28872 12310 28928
rect 14554 31728 14610 31784
rect 12714 30912 12770 30968
rect 12714 28908 12716 28928
rect 12716 28908 12768 28928
rect 12768 28908 12770 28928
rect 12714 28872 12770 28908
rect 12622 27920 12678 27976
rect 12622 27784 12678 27840
rect 12438 27104 12494 27160
rect 11978 25880 12034 25936
rect 12530 26732 12532 26752
rect 12532 26732 12584 26752
rect 12584 26732 12586 26752
rect 12530 26696 12586 26732
rect 13082 29996 13084 30016
rect 13084 29996 13136 30016
rect 13136 29996 13138 30016
rect 13082 29960 13138 29996
rect 13174 29824 13230 29880
rect 12898 28872 12954 28928
rect 13174 28464 13230 28520
rect 13634 30368 13690 30424
rect 13358 28192 13414 28248
rect 12990 27276 12992 27296
rect 12992 27276 13044 27296
rect 13044 27276 13046 27296
rect 12990 27240 13046 27276
rect 12990 27104 13046 27160
rect 12438 26324 12440 26344
rect 12440 26324 12492 26344
rect 12492 26324 12494 26344
rect 12438 26288 12494 26324
rect 13174 27412 13176 27432
rect 13176 27412 13228 27432
rect 13228 27412 13230 27432
rect 13174 27376 13230 27412
rect 13174 26988 13230 27024
rect 13174 26968 13176 26988
rect 13176 26968 13228 26988
rect 13228 26968 13230 26988
rect 12622 25744 12678 25800
rect 12990 26016 13046 26072
rect 13450 27920 13506 27976
rect 13450 27240 13506 27296
rect 14848 31578 14904 31580
rect 14928 31578 14984 31580
rect 15008 31578 15064 31580
rect 15088 31578 15144 31580
rect 14848 31526 14894 31578
rect 14894 31526 14904 31578
rect 14928 31526 14958 31578
rect 14958 31526 14970 31578
rect 14970 31526 14984 31578
rect 15008 31526 15022 31578
rect 15022 31526 15034 31578
rect 15034 31526 15064 31578
rect 15088 31526 15098 31578
rect 15098 31526 15144 31578
rect 14848 31524 14904 31526
rect 14928 31524 14984 31526
rect 15008 31524 15064 31526
rect 15088 31524 15144 31526
rect 14278 30640 14334 30696
rect 14186 29144 14242 29200
rect 14094 28600 14150 28656
rect 15382 30912 15438 30968
rect 14848 30490 14904 30492
rect 14928 30490 14984 30492
rect 15008 30490 15064 30492
rect 15088 30490 15144 30492
rect 14848 30438 14894 30490
rect 14894 30438 14904 30490
rect 14928 30438 14958 30490
rect 14958 30438 14970 30490
rect 14970 30438 14984 30490
rect 15008 30438 15022 30490
rect 15022 30438 15034 30490
rect 15034 30438 15064 30490
rect 15088 30438 15098 30490
rect 15098 30438 15144 30490
rect 14848 30436 14904 30438
rect 14928 30436 14984 30438
rect 15008 30436 15064 30438
rect 15088 30436 15144 30438
rect 14554 30368 14610 30424
rect 15566 30368 15622 30424
rect 14646 29824 14702 29880
rect 14830 29824 14886 29880
rect 15014 29688 15070 29744
rect 15474 29688 15530 29744
rect 14646 29452 14648 29472
rect 14648 29452 14700 29472
rect 14700 29452 14702 29472
rect 14646 29416 14702 29452
rect 14848 29402 14904 29404
rect 14928 29402 14984 29404
rect 15008 29402 15064 29404
rect 15088 29402 15144 29404
rect 14848 29350 14894 29402
rect 14894 29350 14904 29402
rect 14928 29350 14958 29402
rect 14958 29350 14970 29402
rect 14970 29350 14984 29402
rect 15008 29350 15022 29402
rect 15022 29350 15034 29402
rect 15034 29350 15064 29402
rect 15088 29350 15098 29402
rect 15098 29350 15144 29402
rect 14848 29348 14904 29350
rect 14928 29348 14984 29350
rect 15008 29348 15064 29350
rect 15088 29348 15144 29350
rect 13910 28464 13966 28520
rect 13450 26832 13506 26888
rect 13818 27648 13874 27704
rect 13910 27376 13966 27432
rect 13634 26444 13690 26480
rect 13634 26424 13636 26444
rect 13636 26424 13688 26444
rect 13688 26424 13690 26444
rect 14186 27648 14242 27704
rect 14094 26968 14150 27024
rect 15382 29300 15438 29336
rect 15382 29280 15384 29300
rect 15384 29280 15436 29300
rect 15436 29280 15438 29300
rect 14738 29008 14794 29064
rect 14848 28314 14904 28316
rect 14928 28314 14984 28316
rect 15008 28314 15064 28316
rect 15088 28314 15144 28316
rect 14848 28262 14894 28314
rect 14894 28262 14904 28314
rect 14928 28262 14958 28314
rect 14958 28262 14970 28314
rect 14970 28262 14984 28314
rect 15008 28262 15022 28314
rect 15022 28262 15034 28314
rect 15034 28262 15064 28314
rect 15088 28262 15098 28314
rect 15098 28262 15144 28314
rect 14848 28260 14904 28262
rect 14928 28260 14984 28262
rect 15008 28260 15064 28262
rect 15088 28260 15144 28262
rect 15014 28076 15070 28112
rect 15014 28056 15016 28076
rect 15016 28056 15068 28076
rect 15068 28056 15070 28076
rect 14848 27226 14904 27228
rect 14928 27226 14984 27228
rect 15008 27226 15064 27228
rect 15088 27226 15144 27228
rect 14848 27174 14894 27226
rect 14894 27174 14904 27226
rect 14928 27174 14958 27226
rect 14958 27174 14970 27226
rect 14970 27174 14984 27226
rect 15008 27174 15022 27226
rect 15022 27174 15034 27226
rect 15034 27174 15064 27226
rect 15088 27174 15098 27226
rect 15098 27174 15144 27226
rect 14848 27172 14904 27174
rect 14928 27172 14984 27174
rect 15008 27172 15064 27174
rect 15088 27172 15144 27174
rect 15842 29552 15898 29608
rect 15474 27956 15476 27976
rect 15476 27956 15528 27976
rect 15528 27956 15530 27976
rect 15474 27920 15530 27956
rect 14094 26288 14150 26344
rect 14462 26696 14518 26752
rect 14848 26138 14904 26140
rect 14928 26138 14984 26140
rect 15008 26138 15064 26140
rect 15088 26138 15144 26140
rect 14848 26086 14894 26138
rect 14894 26086 14904 26138
rect 14928 26086 14958 26138
rect 14958 26086 14970 26138
rect 14970 26086 14984 26138
rect 15008 26086 15022 26138
rect 15022 26086 15034 26138
rect 15034 26086 15064 26138
rect 15088 26086 15098 26138
rect 15098 26086 15144 26138
rect 14848 26084 14904 26086
rect 14928 26084 14984 26086
rect 15008 26084 15064 26086
rect 15088 26084 15144 26086
rect 16210 29688 16266 29744
rect 16210 29416 16266 29472
rect 15658 27376 15714 27432
rect 15934 27548 15936 27568
rect 15936 27548 15988 27568
rect 15988 27548 15990 27568
rect 15934 27512 15990 27548
rect 15750 26968 15806 27024
rect 16486 30640 16542 30696
rect 16670 31048 16726 31104
rect 17866 31048 17922 31104
rect 16578 30232 16634 30288
rect 16670 29416 16726 29472
rect 16670 29164 16726 29200
rect 16670 29144 16672 29164
rect 16672 29144 16724 29164
rect 16724 29144 16726 29164
rect 16762 28872 16818 28928
rect 17130 29824 17186 29880
rect 17038 29008 17094 29064
rect 16302 26288 16358 26344
rect 16026 25880 16082 25936
rect 14848 25050 14904 25052
rect 14928 25050 14984 25052
rect 15008 25050 15064 25052
rect 15088 25050 15144 25052
rect 14848 24998 14894 25050
rect 14894 24998 14904 25050
rect 14928 24998 14958 25050
rect 14958 24998 14970 25050
rect 14970 24998 14984 25050
rect 15008 24998 15022 25050
rect 15022 24998 15034 25050
rect 15034 24998 15064 25050
rect 15088 24998 15098 25050
rect 15098 24998 15144 25050
rect 14848 24996 14904 24998
rect 14928 24996 14984 24998
rect 15008 24996 15064 24998
rect 15088 24996 15144 24998
rect 17314 29552 17370 29608
rect 17130 27648 17186 27704
rect 17314 26696 17370 26752
rect 14848 23962 14904 23964
rect 14928 23962 14984 23964
rect 15008 23962 15064 23964
rect 15088 23962 15144 23964
rect 14848 23910 14894 23962
rect 14894 23910 14904 23962
rect 14928 23910 14958 23962
rect 14958 23910 14970 23962
rect 14970 23910 14984 23962
rect 15008 23910 15022 23962
rect 15022 23910 15034 23962
rect 15034 23910 15064 23962
rect 15088 23910 15098 23962
rect 15098 23910 15144 23962
rect 14848 23908 14904 23910
rect 14928 23908 14984 23910
rect 15008 23908 15064 23910
rect 15088 23908 15144 23910
rect 11375 23418 11431 23420
rect 11455 23418 11511 23420
rect 11535 23418 11591 23420
rect 11615 23418 11671 23420
rect 11375 23366 11421 23418
rect 11421 23366 11431 23418
rect 11455 23366 11485 23418
rect 11485 23366 11497 23418
rect 11497 23366 11511 23418
rect 11535 23366 11549 23418
rect 11549 23366 11561 23418
rect 11561 23366 11591 23418
rect 11615 23366 11625 23418
rect 11625 23366 11671 23418
rect 11375 23364 11431 23366
rect 11455 23364 11511 23366
rect 11535 23364 11591 23366
rect 11615 23364 11671 23366
rect 7902 22874 7958 22876
rect 7982 22874 8038 22876
rect 8062 22874 8118 22876
rect 8142 22874 8198 22876
rect 7902 22822 7948 22874
rect 7948 22822 7958 22874
rect 7982 22822 8012 22874
rect 8012 22822 8024 22874
rect 8024 22822 8038 22874
rect 8062 22822 8076 22874
rect 8076 22822 8088 22874
rect 8088 22822 8118 22874
rect 8142 22822 8152 22874
rect 8152 22822 8198 22874
rect 7902 22820 7958 22822
rect 7982 22820 8038 22822
rect 8062 22820 8118 22822
rect 8142 22820 8198 22822
rect 14848 22874 14904 22876
rect 14928 22874 14984 22876
rect 15008 22874 15064 22876
rect 15088 22874 15144 22876
rect 14848 22822 14894 22874
rect 14894 22822 14904 22874
rect 14928 22822 14958 22874
rect 14958 22822 14970 22874
rect 14970 22822 14984 22874
rect 15008 22822 15022 22874
rect 15022 22822 15034 22874
rect 15034 22822 15064 22874
rect 15088 22822 15098 22874
rect 15098 22822 15144 22874
rect 14848 22820 14904 22822
rect 14928 22820 14984 22822
rect 15008 22820 15064 22822
rect 15088 22820 15144 22822
rect 4429 22330 4485 22332
rect 4509 22330 4565 22332
rect 4589 22330 4645 22332
rect 4669 22330 4725 22332
rect 4429 22278 4475 22330
rect 4475 22278 4485 22330
rect 4509 22278 4539 22330
rect 4539 22278 4551 22330
rect 4551 22278 4565 22330
rect 4589 22278 4603 22330
rect 4603 22278 4615 22330
rect 4615 22278 4645 22330
rect 4669 22278 4679 22330
rect 4679 22278 4725 22330
rect 4429 22276 4485 22278
rect 4509 22276 4565 22278
rect 4589 22276 4645 22278
rect 4669 22276 4725 22278
rect 11375 22330 11431 22332
rect 11455 22330 11511 22332
rect 11535 22330 11591 22332
rect 11615 22330 11671 22332
rect 11375 22278 11421 22330
rect 11421 22278 11431 22330
rect 11455 22278 11485 22330
rect 11485 22278 11497 22330
rect 11497 22278 11511 22330
rect 11535 22278 11549 22330
rect 11549 22278 11561 22330
rect 11561 22278 11591 22330
rect 11615 22278 11625 22330
rect 11625 22278 11671 22330
rect 11375 22276 11431 22278
rect 11455 22276 11511 22278
rect 11535 22276 11591 22278
rect 11615 22276 11671 22278
rect 1582 22072 1638 22128
rect 7902 21786 7958 21788
rect 7982 21786 8038 21788
rect 8062 21786 8118 21788
rect 8142 21786 8198 21788
rect 7902 21734 7948 21786
rect 7948 21734 7958 21786
rect 7982 21734 8012 21786
rect 8012 21734 8024 21786
rect 8024 21734 8038 21786
rect 8062 21734 8076 21786
rect 8076 21734 8088 21786
rect 8088 21734 8118 21786
rect 8142 21734 8152 21786
rect 8152 21734 8198 21786
rect 7902 21732 7958 21734
rect 7982 21732 8038 21734
rect 8062 21732 8118 21734
rect 8142 21732 8198 21734
rect 14848 21786 14904 21788
rect 14928 21786 14984 21788
rect 15008 21786 15064 21788
rect 15088 21786 15144 21788
rect 14848 21734 14894 21786
rect 14894 21734 14904 21786
rect 14928 21734 14958 21786
rect 14958 21734 14970 21786
rect 14970 21734 14984 21786
rect 15008 21734 15022 21786
rect 15022 21734 15034 21786
rect 15034 21734 15064 21786
rect 15088 21734 15098 21786
rect 15098 21734 15144 21786
rect 14848 21732 14904 21734
rect 14928 21732 14984 21734
rect 15008 21732 15064 21734
rect 15088 21732 15144 21734
rect 1582 21428 1584 21448
rect 1584 21428 1636 21448
rect 1636 21428 1638 21448
rect 1582 21392 1638 21428
rect 4429 21242 4485 21244
rect 4509 21242 4565 21244
rect 4589 21242 4645 21244
rect 4669 21242 4725 21244
rect 4429 21190 4475 21242
rect 4475 21190 4485 21242
rect 4509 21190 4539 21242
rect 4539 21190 4551 21242
rect 4551 21190 4565 21242
rect 4589 21190 4603 21242
rect 4603 21190 4615 21242
rect 4615 21190 4645 21242
rect 4669 21190 4679 21242
rect 4679 21190 4725 21242
rect 4429 21188 4485 21190
rect 4509 21188 4565 21190
rect 4589 21188 4645 21190
rect 4669 21188 4725 21190
rect 11375 21242 11431 21244
rect 11455 21242 11511 21244
rect 11535 21242 11591 21244
rect 11615 21242 11671 21244
rect 11375 21190 11421 21242
rect 11421 21190 11431 21242
rect 11455 21190 11485 21242
rect 11485 21190 11497 21242
rect 11497 21190 11511 21242
rect 11535 21190 11549 21242
rect 11549 21190 11561 21242
rect 11561 21190 11591 21242
rect 11615 21190 11625 21242
rect 11625 21190 11671 21242
rect 11375 21188 11431 21190
rect 11455 21188 11511 21190
rect 11535 21188 11591 21190
rect 11615 21188 11671 21190
rect 7902 20698 7958 20700
rect 7982 20698 8038 20700
rect 8062 20698 8118 20700
rect 8142 20698 8198 20700
rect 7902 20646 7948 20698
rect 7948 20646 7958 20698
rect 7982 20646 8012 20698
rect 8012 20646 8024 20698
rect 8024 20646 8038 20698
rect 8062 20646 8076 20698
rect 8076 20646 8088 20698
rect 8088 20646 8118 20698
rect 8142 20646 8152 20698
rect 8152 20646 8198 20698
rect 7902 20644 7958 20646
rect 7982 20644 8038 20646
rect 8062 20644 8118 20646
rect 8142 20644 8198 20646
rect 14848 20698 14904 20700
rect 14928 20698 14984 20700
rect 15008 20698 15064 20700
rect 15088 20698 15144 20700
rect 14848 20646 14894 20698
rect 14894 20646 14904 20698
rect 14928 20646 14958 20698
rect 14958 20646 14970 20698
rect 14970 20646 14984 20698
rect 15008 20646 15022 20698
rect 15022 20646 15034 20698
rect 15034 20646 15064 20698
rect 15088 20646 15098 20698
rect 15098 20646 15144 20698
rect 14848 20644 14904 20646
rect 14928 20644 14984 20646
rect 15008 20644 15064 20646
rect 15088 20644 15144 20646
rect 4429 20154 4485 20156
rect 4509 20154 4565 20156
rect 4589 20154 4645 20156
rect 4669 20154 4725 20156
rect 4429 20102 4475 20154
rect 4475 20102 4485 20154
rect 4509 20102 4539 20154
rect 4539 20102 4551 20154
rect 4551 20102 4565 20154
rect 4589 20102 4603 20154
rect 4603 20102 4615 20154
rect 4615 20102 4645 20154
rect 4669 20102 4679 20154
rect 4679 20102 4725 20154
rect 4429 20100 4485 20102
rect 4509 20100 4565 20102
rect 4589 20100 4645 20102
rect 4669 20100 4725 20102
rect 11375 20154 11431 20156
rect 11455 20154 11511 20156
rect 11535 20154 11591 20156
rect 11615 20154 11671 20156
rect 11375 20102 11421 20154
rect 11421 20102 11431 20154
rect 11455 20102 11485 20154
rect 11485 20102 11497 20154
rect 11497 20102 11511 20154
rect 11535 20102 11549 20154
rect 11549 20102 11561 20154
rect 11561 20102 11591 20154
rect 11615 20102 11625 20154
rect 11625 20102 11671 20154
rect 11375 20100 11431 20102
rect 11455 20100 11511 20102
rect 11535 20100 11591 20102
rect 11615 20100 11671 20102
rect 1582 20032 1638 20088
rect 7902 19610 7958 19612
rect 7982 19610 8038 19612
rect 8062 19610 8118 19612
rect 8142 19610 8198 19612
rect 7902 19558 7948 19610
rect 7948 19558 7958 19610
rect 7982 19558 8012 19610
rect 8012 19558 8024 19610
rect 8024 19558 8038 19610
rect 8062 19558 8076 19610
rect 8076 19558 8088 19610
rect 8088 19558 8118 19610
rect 8142 19558 8152 19610
rect 8152 19558 8198 19610
rect 7902 19556 7958 19558
rect 7982 19556 8038 19558
rect 8062 19556 8118 19558
rect 8142 19556 8198 19558
rect 14848 19610 14904 19612
rect 14928 19610 14984 19612
rect 15008 19610 15064 19612
rect 15088 19610 15144 19612
rect 14848 19558 14894 19610
rect 14894 19558 14904 19610
rect 14928 19558 14958 19610
rect 14958 19558 14970 19610
rect 14970 19558 14984 19610
rect 15008 19558 15022 19610
rect 15022 19558 15034 19610
rect 15034 19558 15064 19610
rect 15088 19558 15098 19610
rect 15098 19558 15144 19610
rect 14848 19556 14904 19558
rect 14928 19556 14984 19558
rect 15008 19556 15064 19558
rect 15088 19556 15144 19558
rect 1582 19352 1638 19408
rect 4429 19066 4485 19068
rect 4509 19066 4565 19068
rect 4589 19066 4645 19068
rect 4669 19066 4725 19068
rect 4429 19014 4475 19066
rect 4475 19014 4485 19066
rect 4509 19014 4539 19066
rect 4539 19014 4551 19066
rect 4551 19014 4565 19066
rect 4589 19014 4603 19066
rect 4603 19014 4615 19066
rect 4615 19014 4645 19066
rect 4669 19014 4679 19066
rect 4679 19014 4725 19066
rect 4429 19012 4485 19014
rect 4509 19012 4565 19014
rect 4589 19012 4645 19014
rect 4669 19012 4725 19014
rect 11375 19066 11431 19068
rect 11455 19066 11511 19068
rect 11535 19066 11591 19068
rect 11615 19066 11671 19068
rect 11375 19014 11421 19066
rect 11421 19014 11431 19066
rect 11455 19014 11485 19066
rect 11485 19014 11497 19066
rect 11497 19014 11511 19066
rect 11535 19014 11549 19066
rect 11549 19014 11561 19066
rect 11561 19014 11591 19066
rect 11615 19014 11625 19066
rect 11625 19014 11671 19066
rect 11375 19012 11431 19014
rect 11455 19012 11511 19014
rect 11535 19012 11591 19014
rect 11615 19012 11671 19014
rect 7902 18522 7958 18524
rect 7982 18522 8038 18524
rect 8062 18522 8118 18524
rect 8142 18522 8198 18524
rect 7902 18470 7948 18522
rect 7948 18470 7958 18522
rect 7982 18470 8012 18522
rect 8012 18470 8024 18522
rect 8024 18470 8038 18522
rect 8062 18470 8076 18522
rect 8076 18470 8088 18522
rect 8088 18470 8118 18522
rect 8142 18470 8152 18522
rect 8152 18470 8198 18522
rect 7902 18468 7958 18470
rect 7982 18468 8038 18470
rect 8062 18468 8118 18470
rect 8142 18468 8198 18470
rect 14848 18522 14904 18524
rect 14928 18522 14984 18524
rect 15008 18522 15064 18524
rect 15088 18522 15144 18524
rect 14848 18470 14894 18522
rect 14894 18470 14904 18522
rect 14928 18470 14958 18522
rect 14958 18470 14970 18522
rect 14970 18470 14984 18522
rect 15008 18470 15022 18522
rect 15022 18470 15034 18522
rect 15034 18470 15064 18522
rect 15088 18470 15098 18522
rect 15098 18470 15144 18522
rect 14848 18468 14904 18470
rect 14928 18468 14984 18470
rect 15008 18468 15064 18470
rect 15088 18468 15144 18470
rect 1582 18028 1584 18048
rect 1584 18028 1636 18048
rect 1636 18028 1638 18048
rect 1582 17992 1638 18028
rect 4429 17978 4485 17980
rect 4509 17978 4565 17980
rect 4589 17978 4645 17980
rect 4669 17978 4725 17980
rect 4429 17926 4475 17978
rect 4475 17926 4485 17978
rect 4509 17926 4539 17978
rect 4539 17926 4551 17978
rect 4551 17926 4565 17978
rect 4589 17926 4603 17978
rect 4603 17926 4615 17978
rect 4615 17926 4645 17978
rect 4669 17926 4679 17978
rect 4679 17926 4725 17978
rect 4429 17924 4485 17926
rect 4509 17924 4565 17926
rect 4589 17924 4645 17926
rect 4669 17924 4725 17926
rect 11375 17978 11431 17980
rect 11455 17978 11511 17980
rect 11535 17978 11591 17980
rect 11615 17978 11671 17980
rect 11375 17926 11421 17978
rect 11421 17926 11431 17978
rect 11455 17926 11485 17978
rect 11485 17926 11497 17978
rect 11497 17926 11511 17978
rect 11535 17926 11549 17978
rect 11549 17926 11561 17978
rect 11561 17926 11591 17978
rect 11615 17926 11625 17978
rect 11625 17926 11671 17978
rect 11375 17924 11431 17926
rect 11455 17924 11511 17926
rect 11535 17924 11591 17926
rect 11615 17924 11671 17926
rect 7902 17434 7958 17436
rect 7982 17434 8038 17436
rect 8062 17434 8118 17436
rect 8142 17434 8198 17436
rect 7902 17382 7948 17434
rect 7948 17382 7958 17434
rect 7982 17382 8012 17434
rect 8012 17382 8024 17434
rect 8024 17382 8038 17434
rect 8062 17382 8076 17434
rect 8076 17382 8088 17434
rect 8088 17382 8118 17434
rect 8142 17382 8152 17434
rect 8152 17382 8198 17434
rect 7902 17380 7958 17382
rect 7982 17380 8038 17382
rect 8062 17380 8118 17382
rect 8142 17380 8198 17382
rect 14848 17434 14904 17436
rect 14928 17434 14984 17436
rect 15008 17434 15064 17436
rect 15088 17434 15144 17436
rect 14848 17382 14894 17434
rect 14894 17382 14904 17434
rect 14928 17382 14958 17434
rect 14958 17382 14970 17434
rect 14970 17382 14984 17434
rect 15008 17382 15022 17434
rect 15022 17382 15034 17434
rect 15034 17382 15064 17434
rect 15088 17382 15098 17434
rect 15098 17382 15144 17434
rect 14848 17380 14904 17382
rect 14928 17380 14984 17382
rect 15008 17380 15064 17382
rect 15088 17380 15144 17382
rect 1582 17312 1638 17368
rect 4429 16890 4485 16892
rect 4509 16890 4565 16892
rect 4589 16890 4645 16892
rect 4669 16890 4725 16892
rect 4429 16838 4475 16890
rect 4475 16838 4485 16890
rect 4509 16838 4539 16890
rect 4539 16838 4551 16890
rect 4551 16838 4565 16890
rect 4589 16838 4603 16890
rect 4603 16838 4615 16890
rect 4615 16838 4645 16890
rect 4669 16838 4679 16890
rect 4679 16838 4725 16890
rect 4429 16836 4485 16838
rect 4509 16836 4565 16838
rect 4589 16836 4645 16838
rect 4669 16836 4725 16838
rect 11375 16890 11431 16892
rect 11455 16890 11511 16892
rect 11535 16890 11591 16892
rect 11615 16890 11671 16892
rect 11375 16838 11421 16890
rect 11421 16838 11431 16890
rect 11455 16838 11485 16890
rect 11485 16838 11497 16890
rect 11497 16838 11511 16890
rect 11535 16838 11549 16890
rect 11549 16838 11561 16890
rect 11561 16838 11591 16890
rect 11615 16838 11625 16890
rect 11625 16838 11671 16890
rect 11375 16836 11431 16838
rect 11455 16836 11511 16838
rect 11535 16836 11591 16838
rect 11615 16836 11671 16838
rect 7902 16346 7958 16348
rect 7982 16346 8038 16348
rect 8062 16346 8118 16348
rect 8142 16346 8198 16348
rect 7902 16294 7948 16346
rect 7948 16294 7958 16346
rect 7982 16294 8012 16346
rect 8012 16294 8024 16346
rect 8024 16294 8038 16346
rect 8062 16294 8076 16346
rect 8076 16294 8088 16346
rect 8088 16294 8118 16346
rect 8142 16294 8152 16346
rect 8152 16294 8198 16346
rect 7902 16292 7958 16294
rect 7982 16292 8038 16294
rect 8062 16292 8118 16294
rect 8142 16292 8198 16294
rect 14848 16346 14904 16348
rect 14928 16346 14984 16348
rect 15008 16346 15064 16348
rect 15088 16346 15144 16348
rect 14848 16294 14894 16346
rect 14894 16294 14904 16346
rect 14928 16294 14958 16346
rect 14958 16294 14970 16346
rect 14970 16294 14984 16346
rect 15008 16294 15022 16346
rect 15022 16294 15034 16346
rect 15034 16294 15064 16346
rect 15088 16294 15098 16346
rect 15098 16294 15144 16346
rect 14848 16292 14904 16294
rect 14928 16292 14984 16294
rect 15008 16292 15064 16294
rect 15088 16292 15144 16294
rect 1582 15988 1584 16008
rect 1584 15988 1636 16008
rect 1636 15988 1638 16008
rect 1582 15952 1638 15988
rect 4429 15802 4485 15804
rect 4509 15802 4565 15804
rect 4589 15802 4645 15804
rect 4669 15802 4725 15804
rect 4429 15750 4475 15802
rect 4475 15750 4485 15802
rect 4509 15750 4539 15802
rect 4539 15750 4551 15802
rect 4551 15750 4565 15802
rect 4589 15750 4603 15802
rect 4603 15750 4615 15802
rect 4615 15750 4645 15802
rect 4669 15750 4679 15802
rect 4679 15750 4725 15802
rect 4429 15748 4485 15750
rect 4509 15748 4565 15750
rect 4589 15748 4645 15750
rect 4669 15748 4725 15750
rect 11375 15802 11431 15804
rect 11455 15802 11511 15804
rect 11535 15802 11591 15804
rect 11615 15802 11671 15804
rect 11375 15750 11421 15802
rect 11421 15750 11431 15802
rect 11455 15750 11485 15802
rect 11485 15750 11497 15802
rect 11497 15750 11511 15802
rect 11535 15750 11549 15802
rect 11549 15750 11561 15802
rect 11561 15750 11591 15802
rect 11615 15750 11625 15802
rect 11625 15750 11671 15802
rect 11375 15748 11431 15750
rect 11455 15748 11511 15750
rect 11535 15748 11591 15750
rect 11615 15748 11671 15750
rect 1582 15272 1638 15328
rect 7902 15258 7958 15260
rect 7982 15258 8038 15260
rect 8062 15258 8118 15260
rect 8142 15258 8198 15260
rect 7902 15206 7948 15258
rect 7948 15206 7958 15258
rect 7982 15206 8012 15258
rect 8012 15206 8024 15258
rect 8024 15206 8038 15258
rect 8062 15206 8076 15258
rect 8076 15206 8088 15258
rect 8088 15206 8118 15258
rect 8142 15206 8152 15258
rect 8152 15206 8198 15258
rect 7902 15204 7958 15206
rect 7982 15204 8038 15206
rect 8062 15204 8118 15206
rect 8142 15204 8198 15206
rect 14848 15258 14904 15260
rect 14928 15258 14984 15260
rect 15008 15258 15064 15260
rect 15088 15258 15144 15260
rect 14848 15206 14894 15258
rect 14894 15206 14904 15258
rect 14928 15206 14958 15258
rect 14958 15206 14970 15258
rect 14970 15206 14984 15258
rect 15008 15206 15022 15258
rect 15022 15206 15034 15258
rect 15034 15206 15064 15258
rect 15088 15206 15098 15258
rect 15098 15206 15144 15258
rect 14848 15204 14904 15206
rect 14928 15204 14984 15206
rect 15008 15204 15064 15206
rect 15088 15204 15144 15206
rect 4429 14714 4485 14716
rect 4509 14714 4565 14716
rect 4589 14714 4645 14716
rect 4669 14714 4725 14716
rect 4429 14662 4475 14714
rect 4475 14662 4485 14714
rect 4509 14662 4539 14714
rect 4539 14662 4551 14714
rect 4551 14662 4565 14714
rect 4589 14662 4603 14714
rect 4603 14662 4615 14714
rect 4615 14662 4645 14714
rect 4669 14662 4679 14714
rect 4679 14662 4725 14714
rect 4429 14660 4485 14662
rect 4509 14660 4565 14662
rect 4589 14660 4645 14662
rect 4669 14660 4725 14662
rect 11375 14714 11431 14716
rect 11455 14714 11511 14716
rect 11535 14714 11591 14716
rect 11615 14714 11671 14716
rect 11375 14662 11421 14714
rect 11421 14662 11431 14714
rect 11455 14662 11485 14714
rect 11485 14662 11497 14714
rect 11497 14662 11511 14714
rect 11535 14662 11549 14714
rect 11549 14662 11561 14714
rect 11561 14662 11591 14714
rect 11615 14662 11625 14714
rect 11625 14662 11671 14714
rect 11375 14660 11431 14662
rect 11455 14660 11511 14662
rect 11535 14660 11591 14662
rect 11615 14660 11671 14662
rect 7902 14170 7958 14172
rect 7982 14170 8038 14172
rect 8062 14170 8118 14172
rect 8142 14170 8198 14172
rect 7902 14118 7948 14170
rect 7948 14118 7958 14170
rect 7982 14118 8012 14170
rect 8012 14118 8024 14170
rect 8024 14118 8038 14170
rect 8062 14118 8076 14170
rect 8076 14118 8088 14170
rect 8088 14118 8118 14170
rect 8142 14118 8152 14170
rect 8152 14118 8198 14170
rect 7902 14116 7958 14118
rect 7982 14116 8038 14118
rect 8062 14116 8118 14118
rect 8142 14116 8198 14118
rect 14848 14170 14904 14172
rect 14928 14170 14984 14172
rect 15008 14170 15064 14172
rect 15088 14170 15144 14172
rect 14848 14118 14894 14170
rect 14894 14118 14904 14170
rect 14928 14118 14958 14170
rect 14958 14118 14970 14170
rect 14970 14118 14984 14170
rect 15008 14118 15022 14170
rect 15022 14118 15034 14170
rect 15034 14118 15064 14170
rect 15088 14118 15098 14170
rect 15098 14118 15144 14170
rect 14848 14116 14904 14118
rect 14928 14116 14984 14118
rect 15008 14116 15064 14118
rect 15088 14116 15144 14118
rect 1582 13912 1638 13968
rect 4429 13626 4485 13628
rect 4509 13626 4565 13628
rect 4589 13626 4645 13628
rect 4669 13626 4725 13628
rect 4429 13574 4475 13626
rect 4475 13574 4485 13626
rect 4509 13574 4539 13626
rect 4539 13574 4551 13626
rect 4551 13574 4565 13626
rect 4589 13574 4603 13626
rect 4603 13574 4615 13626
rect 4615 13574 4645 13626
rect 4669 13574 4679 13626
rect 4679 13574 4725 13626
rect 4429 13572 4485 13574
rect 4509 13572 4565 13574
rect 4589 13572 4645 13574
rect 4669 13572 4725 13574
rect 11375 13626 11431 13628
rect 11455 13626 11511 13628
rect 11535 13626 11591 13628
rect 11615 13626 11671 13628
rect 11375 13574 11421 13626
rect 11421 13574 11431 13626
rect 11455 13574 11485 13626
rect 11485 13574 11497 13626
rect 11497 13574 11511 13626
rect 11535 13574 11549 13626
rect 11549 13574 11561 13626
rect 11561 13574 11591 13626
rect 11615 13574 11625 13626
rect 11625 13574 11671 13626
rect 11375 13572 11431 13574
rect 11455 13572 11511 13574
rect 11535 13572 11591 13574
rect 11615 13572 11671 13574
rect 1582 13268 1584 13288
rect 1584 13268 1636 13288
rect 1636 13268 1638 13288
rect 1582 13232 1638 13268
rect 7902 13082 7958 13084
rect 7982 13082 8038 13084
rect 8062 13082 8118 13084
rect 8142 13082 8198 13084
rect 7902 13030 7948 13082
rect 7948 13030 7958 13082
rect 7982 13030 8012 13082
rect 8012 13030 8024 13082
rect 8024 13030 8038 13082
rect 8062 13030 8076 13082
rect 8076 13030 8088 13082
rect 8088 13030 8118 13082
rect 8142 13030 8152 13082
rect 8152 13030 8198 13082
rect 7902 13028 7958 13030
rect 7982 13028 8038 13030
rect 8062 13028 8118 13030
rect 8142 13028 8198 13030
rect 14848 13082 14904 13084
rect 14928 13082 14984 13084
rect 15008 13082 15064 13084
rect 15088 13082 15144 13084
rect 14848 13030 14894 13082
rect 14894 13030 14904 13082
rect 14928 13030 14958 13082
rect 14958 13030 14970 13082
rect 14970 13030 14984 13082
rect 15008 13030 15022 13082
rect 15022 13030 15034 13082
rect 15034 13030 15064 13082
rect 15088 13030 15098 13082
rect 15098 13030 15144 13082
rect 14848 13028 14904 13030
rect 14928 13028 14984 13030
rect 15008 13028 15064 13030
rect 15088 13028 15144 13030
rect 4429 12538 4485 12540
rect 4509 12538 4565 12540
rect 4589 12538 4645 12540
rect 4669 12538 4725 12540
rect 4429 12486 4475 12538
rect 4475 12486 4485 12538
rect 4509 12486 4539 12538
rect 4539 12486 4551 12538
rect 4551 12486 4565 12538
rect 4589 12486 4603 12538
rect 4603 12486 4615 12538
rect 4615 12486 4645 12538
rect 4669 12486 4679 12538
rect 4679 12486 4725 12538
rect 4429 12484 4485 12486
rect 4509 12484 4565 12486
rect 4589 12484 4645 12486
rect 4669 12484 4725 12486
rect 11375 12538 11431 12540
rect 11455 12538 11511 12540
rect 11535 12538 11591 12540
rect 11615 12538 11671 12540
rect 11375 12486 11421 12538
rect 11421 12486 11431 12538
rect 11455 12486 11485 12538
rect 11485 12486 11497 12538
rect 11497 12486 11511 12538
rect 11535 12486 11549 12538
rect 11549 12486 11561 12538
rect 11561 12486 11591 12538
rect 11615 12486 11625 12538
rect 11625 12486 11671 12538
rect 11375 12484 11431 12486
rect 11455 12484 11511 12486
rect 11535 12484 11591 12486
rect 11615 12484 11671 12486
rect 7902 11994 7958 11996
rect 7982 11994 8038 11996
rect 8062 11994 8118 11996
rect 8142 11994 8198 11996
rect 7902 11942 7948 11994
rect 7948 11942 7958 11994
rect 7982 11942 8012 11994
rect 8012 11942 8024 11994
rect 8024 11942 8038 11994
rect 8062 11942 8076 11994
rect 8076 11942 8088 11994
rect 8088 11942 8118 11994
rect 8142 11942 8152 11994
rect 8152 11942 8198 11994
rect 7902 11940 7958 11942
rect 7982 11940 8038 11942
rect 8062 11940 8118 11942
rect 8142 11940 8198 11942
rect 14848 11994 14904 11996
rect 14928 11994 14984 11996
rect 15008 11994 15064 11996
rect 15088 11994 15144 11996
rect 14848 11942 14894 11994
rect 14894 11942 14904 11994
rect 14928 11942 14958 11994
rect 14958 11942 14970 11994
rect 14970 11942 14984 11994
rect 15008 11942 15022 11994
rect 15022 11942 15034 11994
rect 15034 11942 15064 11994
rect 15088 11942 15098 11994
rect 15098 11942 15144 11994
rect 14848 11940 14904 11942
rect 14928 11940 14984 11942
rect 15008 11940 15064 11942
rect 15088 11940 15144 11942
rect 1582 11872 1638 11928
rect 4429 11450 4485 11452
rect 4509 11450 4565 11452
rect 4589 11450 4645 11452
rect 4669 11450 4725 11452
rect 4429 11398 4475 11450
rect 4475 11398 4485 11450
rect 4509 11398 4539 11450
rect 4539 11398 4551 11450
rect 4551 11398 4565 11450
rect 4589 11398 4603 11450
rect 4603 11398 4615 11450
rect 4615 11398 4645 11450
rect 4669 11398 4679 11450
rect 4679 11398 4725 11450
rect 4429 11396 4485 11398
rect 4509 11396 4565 11398
rect 4589 11396 4645 11398
rect 4669 11396 4725 11398
rect 11375 11450 11431 11452
rect 11455 11450 11511 11452
rect 11535 11450 11591 11452
rect 11615 11450 11671 11452
rect 11375 11398 11421 11450
rect 11421 11398 11431 11450
rect 11455 11398 11485 11450
rect 11485 11398 11497 11450
rect 11497 11398 11511 11450
rect 11535 11398 11549 11450
rect 11549 11398 11561 11450
rect 11561 11398 11591 11450
rect 11615 11398 11625 11450
rect 11625 11398 11671 11450
rect 11375 11396 11431 11398
rect 11455 11396 11511 11398
rect 11535 11396 11591 11398
rect 11615 11396 11671 11398
rect 1582 11192 1638 11248
rect 7902 10906 7958 10908
rect 7982 10906 8038 10908
rect 8062 10906 8118 10908
rect 8142 10906 8198 10908
rect 7902 10854 7948 10906
rect 7948 10854 7958 10906
rect 7982 10854 8012 10906
rect 8012 10854 8024 10906
rect 8024 10854 8038 10906
rect 8062 10854 8076 10906
rect 8076 10854 8088 10906
rect 8088 10854 8118 10906
rect 8142 10854 8152 10906
rect 8152 10854 8198 10906
rect 7902 10852 7958 10854
rect 7982 10852 8038 10854
rect 8062 10852 8118 10854
rect 8142 10852 8198 10854
rect 14848 10906 14904 10908
rect 14928 10906 14984 10908
rect 15008 10906 15064 10908
rect 15088 10906 15144 10908
rect 14848 10854 14894 10906
rect 14894 10854 14904 10906
rect 14928 10854 14958 10906
rect 14958 10854 14970 10906
rect 14970 10854 14984 10906
rect 15008 10854 15022 10906
rect 15022 10854 15034 10906
rect 15034 10854 15064 10906
rect 15088 10854 15098 10906
rect 15098 10854 15144 10906
rect 14848 10852 14904 10854
rect 14928 10852 14984 10854
rect 15008 10852 15064 10854
rect 15088 10852 15144 10854
rect 4429 10362 4485 10364
rect 4509 10362 4565 10364
rect 4589 10362 4645 10364
rect 4669 10362 4725 10364
rect 4429 10310 4475 10362
rect 4475 10310 4485 10362
rect 4509 10310 4539 10362
rect 4539 10310 4551 10362
rect 4551 10310 4565 10362
rect 4589 10310 4603 10362
rect 4603 10310 4615 10362
rect 4615 10310 4645 10362
rect 4669 10310 4679 10362
rect 4679 10310 4725 10362
rect 4429 10308 4485 10310
rect 4509 10308 4565 10310
rect 4589 10308 4645 10310
rect 4669 10308 4725 10310
rect 11375 10362 11431 10364
rect 11455 10362 11511 10364
rect 11535 10362 11591 10364
rect 11615 10362 11671 10364
rect 11375 10310 11421 10362
rect 11421 10310 11431 10362
rect 11455 10310 11485 10362
rect 11485 10310 11497 10362
rect 11497 10310 11511 10362
rect 11535 10310 11549 10362
rect 11549 10310 11561 10362
rect 11561 10310 11591 10362
rect 11615 10310 11625 10362
rect 11625 10310 11671 10362
rect 11375 10308 11431 10310
rect 11455 10308 11511 10310
rect 11535 10308 11591 10310
rect 11615 10308 11671 10310
rect 1582 9832 1638 9888
rect 7902 9818 7958 9820
rect 7982 9818 8038 9820
rect 8062 9818 8118 9820
rect 8142 9818 8198 9820
rect 7902 9766 7948 9818
rect 7948 9766 7958 9818
rect 7982 9766 8012 9818
rect 8012 9766 8024 9818
rect 8024 9766 8038 9818
rect 8062 9766 8076 9818
rect 8076 9766 8088 9818
rect 8088 9766 8118 9818
rect 8142 9766 8152 9818
rect 8152 9766 8198 9818
rect 7902 9764 7958 9766
rect 7982 9764 8038 9766
rect 8062 9764 8118 9766
rect 8142 9764 8198 9766
rect 14848 9818 14904 9820
rect 14928 9818 14984 9820
rect 15008 9818 15064 9820
rect 15088 9818 15144 9820
rect 14848 9766 14894 9818
rect 14894 9766 14904 9818
rect 14928 9766 14958 9818
rect 14958 9766 14970 9818
rect 14970 9766 14984 9818
rect 15008 9766 15022 9818
rect 15022 9766 15034 9818
rect 15034 9766 15064 9818
rect 15088 9766 15098 9818
rect 15098 9766 15144 9818
rect 14848 9764 14904 9766
rect 14928 9764 14984 9766
rect 15008 9764 15064 9766
rect 15088 9764 15144 9766
rect 4429 9274 4485 9276
rect 4509 9274 4565 9276
rect 4589 9274 4645 9276
rect 4669 9274 4725 9276
rect 4429 9222 4475 9274
rect 4475 9222 4485 9274
rect 4509 9222 4539 9274
rect 4539 9222 4551 9274
rect 4551 9222 4565 9274
rect 4589 9222 4603 9274
rect 4603 9222 4615 9274
rect 4615 9222 4645 9274
rect 4669 9222 4679 9274
rect 4679 9222 4725 9274
rect 4429 9220 4485 9222
rect 4509 9220 4565 9222
rect 4589 9220 4645 9222
rect 4669 9220 4725 9222
rect 11375 9274 11431 9276
rect 11455 9274 11511 9276
rect 11535 9274 11591 9276
rect 11615 9274 11671 9276
rect 11375 9222 11421 9274
rect 11421 9222 11431 9274
rect 11455 9222 11485 9274
rect 11485 9222 11497 9274
rect 11497 9222 11511 9274
rect 11535 9222 11549 9274
rect 11549 9222 11561 9274
rect 11561 9222 11591 9274
rect 11615 9222 11625 9274
rect 11625 9222 11671 9274
rect 11375 9220 11431 9222
rect 11455 9220 11511 9222
rect 11535 9220 11591 9222
rect 11615 9220 11671 9222
rect 1582 9152 1638 9208
rect 7902 8730 7958 8732
rect 7982 8730 8038 8732
rect 8062 8730 8118 8732
rect 8142 8730 8198 8732
rect 7902 8678 7948 8730
rect 7948 8678 7958 8730
rect 7982 8678 8012 8730
rect 8012 8678 8024 8730
rect 8024 8678 8038 8730
rect 8062 8678 8076 8730
rect 8076 8678 8088 8730
rect 8088 8678 8118 8730
rect 8142 8678 8152 8730
rect 8152 8678 8198 8730
rect 7902 8676 7958 8678
rect 7982 8676 8038 8678
rect 8062 8676 8118 8678
rect 8142 8676 8198 8678
rect 14848 8730 14904 8732
rect 14928 8730 14984 8732
rect 15008 8730 15064 8732
rect 15088 8730 15144 8732
rect 14848 8678 14894 8730
rect 14894 8678 14904 8730
rect 14928 8678 14958 8730
rect 14958 8678 14970 8730
rect 14970 8678 14984 8730
rect 15008 8678 15022 8730
rect 15022 8678 15034 8730
rect 15034 8678 15064 8730
rect 15088 8678 15098 8730
rect 15098 8678 15144 8730
rect 14848 8676 14904 8678
rect 14928 8676 14984 8678
rect 15008 8676 15064 8678
rect 15088 8676 15144 8678
rect 4429 8186 4485 8188
rect 4509 8186 4565 8188
rect 4589 8186 4645 8188
rect 4669 8186 4725 8188
rect 4429 8134 4475 8186
rect 4475 8134 4485 8186
rect 4509 8134 4539 8186
rect 4539 8134 4551 8186
rect 4551 8134 4565 8186
rect 4589 8134 4603 8186
rect 4603 8134 4615 8186
rect 4615 8134 4645 8186
rect 4669 8134 4679 8186
rect 4679 8134 4725 8186
rect 4429 8132 4485 8134
rect 4509 8132 4565 8134
rect 4589 8132 4645 8134
rect 4669 8132 4725 8134
rect 11375 8186 11431 8188
rect 11455 8186 11511 8188
rect 11535 8186 11591 8188
rect 11615 8186 11671 8188
rect 11375 8134 11421 8186
rect 11421 8134 11431 8186
rect 11455 8134 11485 8186
rect 11485 8134 11497 8186
rect 11497 8134 11511 8186
rect 11535 8134 11549 8186
rect 11549 8134 11561 8186
rect 11561 8134 11591 8186
rect 11615 8134 11625 8186
rect 11625 8134 11671 8186
rect 11375 8132 11431 8134
rect 11455 8132 11511 8134
rect 11535 8132 11591 8134
rect 11615 8132 11671 8134
rect 1582 7828 1584 7848
rect 1584 7828 1636 7848
rect 1636 7828 1638 7848
rect 1582 7792 1638 7828
rect 7902 7642 7958 7644
rect 7982 7642 8038 7644
rect 8062 7642 8118 7644
rect 8142 7642 8198 7644
rect 7902 7590 7948 7642
rect 7948 7590 7958 7642
rect 7982 7590 8012 7642
rect 8012 7590 8024 7642
rect 8024 7590 8038 7642
rect 8062 7590 8076 7642
rect 8076 7590 8088 7642
rect 8088 7590 8118 7642
rect 8142 7590 8152 7642
rect 8152 7590 8198 7642
rect 7902 7588 7958 7590
rect 7982 7588 8038 7590
rect 8062 7588 8118 7590
rect 8142 7588 8198 7590
rect 14848 7642 14904 7644
rect 14928 7642 14984 7644
rect 15008 7642 15064 7644
rect 15088 7642 15144 7644
rect 14848 7590 14894 7642
rect 14894 7590 14904 7642
rect 14928 7590 14958 7642
rect 14958 7590 14970 7642
rect 14970 7590 14984 7642
rect 15008 7590 15022 7642
rect 15022 7590 15034 7642
rect 15034 7590 15064 7642
rect 15088 7590 15098 7642
rect 15098 7590 15144 7642
rect 14848 7588 14904 7590
rect 14928 7588 14984 7590
rect 15008 7588 15064 7590
rect 15088 7588 15144 7590
rect 1582 7148 1584 7168
rect 1584 7148 1636 7168
rect 1636 7148 1638 7168
rect 1582 7112 1638 7148
rect 4429 7098 4485 7100
rect 4509 7098 4565 7100
rect 4589 7098 4645 7100
rect 4669 7098 4725 7100
rect 4429 7046 4475 7098
rect 4475 7046 4485 7098
rect 4509 7046 4539 7098
rect 4539 7046 4551 7098
rect 4551 7046 4565 7098
rect 4589 7046 4603 7098
rect 4603 7046 4615 7098
rect 4615 7046 4645 7098
rect 4669 7046 4679 7098
rect 4679 7046 4725 7098
rect 4429 7044 4485 7046
rect 4509 7044 4565 7046
rect 4589 7044 4645 7046
rect 4669 7044 4725 7046
rect 11375 7098 11431 7100
rect 11455 7098 11511 7100
rect 11535 7098 11591 7100
rect 11615 7098 11671 7100
rect 11375 7046 11421 7098
rect 11421 7046 11431 7098
rect 11455 7046 11485 7098
rect 11485 7046 11497 7098
rect 11497 7046 11511 7098
rect 11535 7046 11549 7098
rect 11549 7046 11561 7098
rect 11561 7046 11591 7098
rect 11615 7046 11625 7098
rect 11625 7046 11671 7098
rect 11375 7044 11431 7046
rect 11455 7044 11511 7046
rect 11535 7044 11591 7046
rect 11615 7044 11671 7046
rect 7902 6554 7958 6556
rect 7982 6554 8038 6556
rect 8062 6554 8118 6556
rect 8142 6554 8198 6556
rect 7902 6502 7948 6554
rect 7948 6502 7958 6554
rect 7982 6502 8012 6554
rect 8012 6502 8024 6554
rect 8024 6502 8038 6554
rect 8062 6502 8076 6554
rect 8076 6502 8088 6554
rect 8088 6502 8118 6554
rect 8142 6502 8152 6554
rect 8152 6502 8198 6554
rect 7902 6500 7958 6502
rect 7982 6500 8038 6502
rect 8062 6500 8118 6502
rect 8142 6500 8198 6502
rect 14848 6554 14904 6556
rect 14928 6554 14984 6556
rect 15008 6554 15064 6556
rect 15088 6554 15144 6556
rect 14848 6502 14894 6554
rect 14894 6502 14904 6554
rect 14928 6502 14958 6554
rect 14958 6502 14970 6554
rect 14970 6502 14984 6554
rect 15008 6502 15022 6554
rect 15022 6502 15034 6554
rect 15034 6502 15064 6554
rect 15088 6502 15098 6554
rect 15098 6502 15144 6554
rect 14848 6500 14904 6502
rect 14928 6500 14984 6502
rect 15008 6500 15064 6502
rect 15088 6500 15144 6502
rect 4429 6010 4485 6012
rect 4509 6010 4565 6012
rect 4589 6010 4645 6012
rect 4669 6010 4725 6012
rect 4429 5958 4475 6010
rect 4475 5958 4485 6010
rect 4509 5958 4539 6010
rect 4539 5958 4551 6010
rect 4551 5958 4565 6010
rect 4589 5958 4603 6010
rect 4603 5958 4615 6010
rect 4615 5958 4645 6010
rect 4669 5958 4679 6010
rect 4679 5958 4725 6010
rect 4429 5956 4485 5958
rect 4509 5956 4565 5958
rect 4589 5956 4645 5958
rect 4669 5956 4725 5958
rect 11375 6010 11431 6012
rect 11455 6010 11511 6012
rect 11535 6010 11591 6012
rect 11615 6010 11671 6012
rect 11375 5958 11421 6010
rect 11421 5958 11431 6010
rect 11455 5958 11485 6010
rect 11485 5958 11497 6010
rect 11497 5958 11511 6010
rect 11535 5958 11549 6010
rect 11549 5958 11561 6010
rect 11561 5958 11591 6010
rect 11615 5958 11625 6010
rect 11625 5958 11671 6010
rect 11375 5956 11431 5958
rect 11455 5956 11511 5958
rect 11535 5956 11591 5958
rect 11615 5956 11671 5958
rect 1582 5752 1638 5808
rect 7902 5466 7958 5468
rect 7982 5466 8038 5468
rect 8062 5466 8118 5468
rect 8142 5466 8198 5468
rect 7902 5414 7948 5466
rect 7948 5414 7958 5466
rect 7982 5414 8012 5466
rect 8012 5414 8024 5466
rect 8024 5414 8038 5466
rect 8062 5414 8076 5466
rect 8076 5414 8088 5466
rect 8088 5414 8118 5466
rect 8142 5414 8152 5466
rect 8152 5414 8198 5466
rect 7902 5412 7958 5414
rect 7982 5412 8038 5414
rect 8062 5412 8118 5414
rect 8142 5412 8198 5414
rect 14848 5466 14904 5468
rect 14928 5466 14984 5468
rect 15008 5466 15064 5468
rect 15088 5466 15144 5468
rect 14848 5414 14894 5466
rect 14894 5414 14904 5466
rect 14928 5414 14958 5466
rect 14958 5414 14970 5466
rect 14970 5414 14984 5466
rect 15008 5414 15022 5466
rect 15022 5414 15034 5466
rect 15034 5414 15064 5466
rect 15088 5414 15098 5466
rect 15098 5414 15144 5466
rect 14848 5412 14904 5414
rect 14928 5412 14984 5414
rect 15008 5412 15064 5414
rect 15088 5412 15144 5414
rect 1582 5108 1584 5128
rect 1584 5108 1636 5128
rect 1636 5108 1638 5128
rect 1582 5072 1638 5108
rect 4429 4922 4485 4924
rect 4509 4922 4565 4924
rect 4589 4922 4645 4924
rect 4669 4922 4725 4924
rect 4429 4870 4475 4922
rect 4475 4870 4485 4922
rect 4509 4870 4539 4922
rect 4539 4870 4551 4922
rect 4551 4870 4565 4922
rect 4589 4870 4603 4922
rect 4603 4870 4615 4922
rect 4615 4870 4645 4922
rect 4669 4870 4679 4922
rect 4679 4870 4725 4922
rect 4429 4868 4485 4870
rect 4509 4868 4565 4870
rect 4589 4868 4645 4870
rect 4669 4868 4725 4870
rect 11375 4922 11431 4924
rect 11455 4922 11511 4924
rect 11535 4922 11591 4924
rect 11615 4922 11671 4924
rect 11375 4870 11421 4922
rect 11421 4870 11431 4922
rect 11455 4870 11485 4922
rect 11485 4870 11497 4922
rect 11497 4870 11511 4922
rect 11535 4870 11549 4922
rect 11549 4870 11561 4922
rect 11561 4870 11591 4922
rect 11615 4870 11625 4922
rect 11625 4870 11671 4922
rect 11375 4868 11431 4870
rect 11455 4868 11511 4870
rect 11535 4868 11591 4870
rect 11615 4868 11671 4870
rect 7902 4378 7958 4380
rect 7982 4378 8038 4380
rect 8062 4378 8118 4380
rect 8142 4378 8198 4380
rect 7902 4326 7948 4378
rect 7948 4326 7958 4378
rect 7982 4326 8012 4378
rect 8012 4326 8024 4378
rect 8024 4326 8038 4378
rect 8062 4326 8076 4378
rect 8076 4326 8088 4378
rect 8088 4326 8118 4378
rect 8142 4326 8152 4378
rect 8152 4326 8198 4378
rect 7902 4324 7958 4326
rect 7982 4324 8038 4326
rect 8062 4324 8118 4326
rect 8142 4324 8198 4326
rect 14848 4378 14904 4380
rect 14928 4378 14984 4380
rect 15008 4378 15064 4380
rect 15088 4378 15144 4380
rect 14848 4326 14894 4378
rect 14894 4326 14904 4378
rect 14928 4326 14958 4378
rect 14958 4326 14970 4378
rect 14970 4326 14984 4378
rect 15008 4326 15022 4378
rect 15022 4326 15034 4378
rect 15034 4326 15064 4378
rect 15088 4326 15098 4378
rect 15098 4326 15144 4378
rect 14848 4324 14904 4326
rect 14928 4324 14984 4326
rect 15008 4324 15064 4326
rect 15088 4324 15144 4326
rect 17498 26560 17554 26616
rect 18694 31184 18750 31240
rect 18321 31034 18377 31036
rect 18401 31034 18457 31036
rect 18481 31034 18537 31036
rect 18561 31034 18617 31036
rect 18321 30982 18367 31034
rect 18367 30982 18377 31034
rect 18401 30982 18431 31034
rect 18431 30982 18443 31034
rect 18443 30982 18457 31034
rect 18481 30982 18495 31034
rect 18495 30982 18507 31034
rect 18507 30982 18537 31034
rect 18561 30982 18571 31034
rect 18571 30982 18617 31034
rect 18321 30980 18377 30982
rect 18401 30980 18457 30982
rect 18481 30980 18537 30982
rect 18561 30980 18617 30982
rect 18321 29946 18377 29948
rect 18401 29946 18457 29948
rect 18481 29946 18537 29948
rect 18561 29946 18617 29948
rect 18321 29894 18367 29946
rect 18367 29894 18377 29946
rect 18401 29894 18431 29946
rect 18431 29894 18443 29946
rect 18443 29894 18457 29946
rect 18481 29894 18495 29946
rect 18495 29894 18507 29946
rect 18507 29894 18537 29946
rect 18561 29894 18571 29946
rect 18571 29894 18617 29946
rect 18321 29892 18377 29894
rect 18401 29892 18457 29894
rect 18481 29892 18537 29894
rect 18561 29892 18617 29894
rect 18142 28736 18198 28792
rect 17958 27784 18014 27840
rect 18321 28858 18377 28860
rect 18401 28858 18457 28860
rect 18481 28858 18537 28860
rect 18561 28858 18617 28860
rect 18321 28806 18367 28858
rect 18367 28806 18377 28858
rect 18401 28806 18431 28858
rect 18431 28806 18443 28858
rect 18443 28806 18457 28858
rect 18481 28806 18495 28858
rect 18495 28806 18507 28858
rect 18507 28806 18537 28858
rect 18561 28806 18571 28858
rect 18571 28806 18617 28858
rect 18321 28804 18377 28806
rect 18401 28804 18457 28806
rect 18481 28804 18537 28806
rect 18561 28804 18617 28806
rect 18970 29552 19026 29608
rect 19798 30812 19800 30832
rect 19800 30812 19852 30832
rect 19852 30812 19854 30832
rect 19798 30776 19854 30812
rect 19890 30368 19946 30424
rect 19614 30096 19670 30152
rect 21794 31578 21850 31580
rect 21874 31578 21930 31580
rect 21954 31578 22010 31580
rect 22034 31578 22090 31580
rect 21794 31526 21840 31578
rect 21840 31526 21850 31578
rect 21874 31526 21904 31578
rect 21904 31526 21916 31578
rect 21916 31526 21930 31578
rect 21954 31526 21968 31578
rect 21968 31526 21980 31578
rect 21980 31526 22010 31578
rect 22034 31526 22044 31578
rect 22044 31526 22090 31578
rect 21794 31524 21850 31526
rect 21874 31524 21930 31526
rect 21954 31524 22010 31526
rect 22034 31524 22090 31526
rect 27710 31864 27766 31920
rect 25267 31034 25323 31036
rect 25347 31034 25403 31036
rect 25427 31034 25483 31036
rect 25507 31034 25563 31036
rect 25267 30982 25313 31034
rect 25313 30982 25323 31034
rect 25347 30982 25377 31034
rect 25377 30982 25389 31034
rect 25389 30982 25403 31034
rect 25427 30982 25441 31034
rect 25441 30982 25453 31034
rect 25453 30982 25483 31034
rect 25507 30982 25517 31034
rect 25517 30982 25563 31034
rect 25267 30980 25323 30982
rect 25347 30980 25403 30982
rect 25427 30980 25483 30982
rect 25507 30980 25563 30982
rect 28740 31578 28796 31580
rect 28820 31578 28876 31580
rect 28900 31578 28956 31580
rect 28980 31578 29036 31580
rect 28740 31526 28786 31578
rect 28786 31526 28796 31578
rect 28820 31526 28850 31578
rect 28850 31526 28862 31578
rect 28862 31526 28876 31578
rect 28900 31526 28914 31578
rect 28914 31526 28926 31578
rect 28926 31526 28956 31578
rect 28980 31526 28990 31578
rect 28990 31526 29036 31578
rect 28740 31524 28796 31526
rect 28820 31524 28876 31526
rect 28900 31524 28956 31526
rect 28980 31524 29036 31526
rect 28354 31184 28410 31240
rect 21794 30490 21850 30492
rect 21874 30490 21930 30492
rect 21954 30490 22010 30492
rect 22034 30490 22090 30492
rect 21794 30438 21840 30490
rect 21840 30438 21850 30490
rect 21874 30438 21904 30490
rect 21904 30438 21916 30490
rect 21916 30438 21930 30490
rect 21954 30438 21968 30490
rect 21968 30438 21980 30490
rect 21980 30438 22010 30490
rect 22034 30438 22044 30490
rect 22044 30438 22090 30490
rect 21794 30436 21850 30438
rect 21874 30436 21930 30438
rect 21954 30436 22010 30438
rect 22034 30436 22090 30438
rect 28740 30490 28796 30492
rect 28820 30490 28876 30492
rect 28900 30490 28956 30492
rect 28980 30490 29036 30492
rect 28740 30438 28786 30490
rect 28786 30438 28796 30490
rect 28820 30438 28850 30490
rect 28850 30438 28862 30490
rect 28862 30438 28876 30490
rect 28900 30438 28914 30490
rect 28914 30438 28926 30490
rect 28926 30438 28956 30490
rect 28980 30438 28990 30490
rect 28990 30438 29036 30490
rect 28740 30436 28796 30438
rect 28820 30436 28876 30438
rect 28900 30436 28956 30438
rect 28980 30436 29036 30438
rect 25267 29946 25323 29948
rect 25347 29946 25403 29948
rect 25427 29946 25483 29948
rect 25507 29946 25563 29948
rect 25267 29894 25313 29946
rect 25313 29894 25323 29946
rect 25347 29894 25377 29946
rect 25377 29894 25389 29946
rect 25389 29894 25403 29946
rect 25427 29894 25441 29946
rect 25441 29894 25453 29946
rect 25453 29894 25483 29946
rect 25507 29894 25517 29946
rect 25517 29894 25563 29946
rect 25267 29892 25323 29894
rect 25347 29892 25403 29894
rect 25427 29892 25483 29894
rect 25507 29892 25563 29894
rect 28354 29824 28410 29880
rect 21794 29402 21850 29404
rect 21874 29402 21930 29404
rect 21954 29402 22010 29404
rect 22034 29402 22090 29404
rect 21794 29350 21840 29402
rect 21840 29350 21850 29402
rect 21874 29350 21904 29402
rect 21904 29350 21916 29402
rect 21916 29350 21930 29402
rect 21954 29350 21968 29402
rect 21968 29350 21980 29402
rect 21980 29350 22010 29402
rect 22034 29350 22044 29402
rect 22044 29350 22090 29402
rect 21794 29348 21850 29350
rect 21874 29348 21930 29350
rect 21954 29348 22010 29350
rect 22034 29348 22090 29350
rect 19062 29280 19118 29336
rect 28740 29402 28796 29404
rect 28820 29402 28876 29404
rect 28900 29402 28956 29404
rect 28980 29402 29036 29404
rect 28740 29350 28786 29402
rect 28786 29350 28796 29402
rect 28820 29350 28850 29402
rect 28850 29350 28862 29402
rect 28862 29350 28876 29402
rect 28900 29350 28914 29402
rect 28914 29350 28926 29402
rect 28926 29350 28956 29402
rect 28980 29350 28990 29402
rect 28990 29350 29036 29402
rect 28740 29348 28796 29350
rect 28820 29348 28876 29350
rect 28900 29348 28956 29350
rect 28980 29348 29036 29350
rect 28354 29144 28410 29200
rect 25267 28858 25323 28860
rect 25347 28858 25403 28860
rect 25427 28858 25483 28860
rect 25507 28858 25563 28860
rect 25267 28806 25313 28858
rect 25313 28806 25323 28858
rect 25347 28806 25377 28858
rect 25377 28806 25389 28858
rect 25389 28806 25403 28858
rect 25427 28806 25441 28858
rect 25441 28806 25453 28858
rect 25453 28806 25483 28858
rect 25507 28806 25517 28858
rect 25517 28806 25563 28858
rect 25267 28804 25323 28806
rect 25347 28804 25403 28806
rect 25427 28804 25483 28806
rect 25507 28804 25563 28806
rect 21794 28314 21850 28316
rect 21874 28314 21930 28316
rect 21954 28314 22010 28316
rect 22034 28314 22090 28316
rect 21794 28262 21840 28314
rect 21840 28262 21850 28314
rect 21874 28262 21904 28314
rect 21904 28262 21916 28314
rect 21916 28262 21930 28314
rect 21954 28262 21968 28314
rect 21968 28262 21980 28314
rect 21980 28262 22010 28314
rect 22034 28262 22044 28314
rect 22044 28262 22090 28314
rect 21794 28260 21850 28262
rect 21874 28260 21930 28262
rect 21954 28260 22010 28262
rect 22034 28260 22090 28262
rect 28740 28314 28796 28316
rect 28820 28314 28876 28316
rect 28900 28314 28956 28316
rect 28980 28314 29036 28316
rect 28740 28262 28786 28314
rect 28786 28262 28796 28314
rect 28820 28262 28850 28314
rect 28850 28262 28862 28314
rect 28862 28262 28876 28314
rect 28900 28262 28914 28314
rect 28914 28262 28926 28314
rect 28926 28262 28956 28314
rect 28980 28262 28990 28314
rect 28990 28262 29036 28314
rect 28740 28260 28796 28262
rect 28820 28260 28876 28262
rect 28900 28260 28956 28262
rect 28980 28260 29036 28262
rect 28354 27820 28356 27840
rect 28356 27820 28408 27840
rect 28408 27820 28410 27840
rect 28354 27784 28410 27820
rect 18321 27770 18377 27772
rect 18401 27770 18457 27772
rect 18481 27770 18537 27772
rect 18561 27770 18617 27772
rect 18321 27718 18367 27770
rect 18367 27718 18377 27770
rect 18401 27718 18431 27770
rect 18431 27718 18443 27770
rect 18443 27718 18457 27770
rect 18481 27718 18495 27770
rect 18495 27718 18507 27770
rect 18507 27718 18537 27770
rect 18561 27718 18571 27770
rect 18571 27718 18617 27770
rect 18321 27716 18377 27718
rect 18401 27716 18457 27718
rect 18481 27716 18537 27718
rect 18561 27716 18617 27718
rect 25267 27770 25323 27772
rect 25347 27770 25403 27772
rect 25427 27770 25483 27772
rect 25507 27770 25563 27772
rect 25267 27718 25313 27770
rect 25313 27718 25323 27770
rect 25347 27718 25377 27770
rect 25377 27718 25389 27770
rect 25389 27718 25403 27770
rect 25427 27718 25441 27770
rect 25441 27718 25453 27770
rect 25453 27718 25483 27770
rect 25507 27718 25517 27770
rect 25517 27718 25563 27770
rect 25267 27716 25323 27718
rect 25347 27716 25403 27718
rect 25427 27716 25483 27718
rect 25507 27716 25563 27718
rect 28354 27412 28356 27432
rect 28356 27412 28408 27432
rect 28408 27412 28410 27432
rect 28354 27376 28410 27412
rect 21794 27226 21850 27228
rect 21874 27226 21930 27228
rect 21954 27226 22010 27228
rect 22034 27226 22090 27228
rect 21794 27174 21840 27226
rect 21840 27174 21850 27226
rect 21874 27174 21904 27226
rect 21904 27174 21916 27226
rect 21916 27174 21930 27226
rect 21954 27174 21968 27226
rect 21968 27174 21980 27226
rect 21980 27174 22010 27226
rect 22034 27174 22044 27226
rect 22044 27174 22090 27226
rect 21794 27172 21850 27174
rect 21874 27172 21930 27174
rect 21954 27172 22010 27174
rect 22034 27172 22090 27174
rect 28740 27226 28796 27228
rect 28820 27226 28876 27228
rect 28900 27226 28956 27228
rect 28980 27226 29036 27228
rect 28740 27174 28786 27226
rect 28786 27174 28796 27226
rect 28820 27174 28850 27226
rect 28850 27174 28862 27226
rect 28862 27174 28876 27226
rect 28900 27174 28914 27226
rect 28914 27174 28926 27226
rect 28926 27174 28956 27226
rect 28980 27174 28990 27226
rect 28990 27174 29036 27226
rect 28740 27172 28796 27174
rect 28820 27172 28876 27174
rect 28900 27172 28956 27174
rect 28980 27172 29036 27174
rect 18321 26682 18377 26684
rect 18401 26682 18457 26684
rect 18481 26682 18537 26684
rect 18561 26682 18617 26684
rect 18321 26630 18367 26682
rect 18367 26630 18377 26682
rect 18401 26630 18431 26682
rect 18431 26630 18443 26682
rect 18443 26630 18457 26682
rect 18481 26630 18495 26682
rect 18495 26630 18507 26682
rect 18507 26630 18537 26682
rect 18561 26630 18571 26682
rect 18571 26630 18617 26682
rect 18321 26628 18377 26630
rect 18401 26628 18457 26630
rect 18481 26628 18537 26630
rect 18561 26628 18617 26630
rect 25267 26682 25323 26684
rect 25347 26682 25403 26684
rect 25427 26682 25483 26684
rect 25507 26682 25563 26684
rect 25267 26630 25313 26682
rect 25313 26630 25323 26682
rect 25347 26630 25377 26682
rect 25377 26630 25389 26682
rect 25389 26630 25403 26682
rect 25427 26630 25441 26682
rect 25441 26630 25453 26682
rect 25453 26630 25483 26682
rect 25507 26630 25517 26682
rect 25517 26630 25563 26682
rect 25267 26628 25323 26630
rect 25347 26628 25403 26630
rect 25427 26628 25483 26630
rect 25507 26628 25563 26630
rect 21794 26138 21850 26140
rect 21874 26138 21930 26140
rect 21954 26138 22010 26140
rect 22034 26138 22090 26140
rect 21794 26086 21840 26138
rect 21840 26086 21850 26138
rect 21874 26086 21904 26138
rect 21904 26086 21916 26138
rect 21916 26086 21930 26138
rect 21954 26086 21968 26138
rect 21968 26086 21980 26138
rect 21980 26086 22010 26138
rect 22034 26086 22044 26138
rect 22044 26086 22090 26138
rect 21794 26084 21850 26086
rect 21874 26084 21930 26086
rect 21954 26084 22010 26086
rect 22034 26084 22090 26086
rect 28740 26138 28796 26140
rect 28820 26138 28876 26140
rect 28900 26138 28956 26140
rect 28980 26138 29036 26140
rect 28740 26086 28786 26138
rect 28786 26086 28796 26138
rect 28820 26086 28850 26138
rect 28850 26086 28862 26138
rect 28862 26086 28876 26138
rect 28900 26086 28914 26138
rect 28914 26086 28926 26138
rect 28926 26086 28956 26138
rect 28980 26086 28990 26138
rect 28990 26086 29036 26138
rect 28740 26084 28796 26086
rect 28820 26084 28876 26086
rect 28900 26084 28956 26086
rect 28980 26084 29036 26086
rect 28354 25764 28410 25800
rect 28354 25744 28356 25764
rect 28356 25744 28408 25764
rect 28408 25744 28410 25764
rect 18321 25594 18377 25596
rect 18401 25594 18457 25596
rect 18481 25594 18537 25596
rect 18561 25594 18617 25596
rect 18321 25542 18367 25594
rect 18367 25542 18377 25594
rect 18401 25542 18431 25594
rect 18431 25542 18443 25594
rect 18443 25542 18457 25594
rect 18481 25542 18495 25594
rect 18495 25542 18507 25594
rect 18507 25542 18537 25594
rect 18561 25542 18571 25594
rect 18571 25542 18617 25594
rect 18321 25540 18377 25542
rect 18401 25540 18457 25542
rect 18481 25540 18537 25542
rect 18561 25540 18617 25542
rect 25267 25594 25323 25596
rect 25347 25594 25403 25596
rect 25427 25594 25483 25596
rect 25507 25594 25563 25596
rect 25267 25542 25313 25594
rect 25313 25542 25323 25594
rect 25347 25542 25377 25594
rect 25377 25542 25389 25594
rect 25389 25542 25403 25594
rect 25427 25542 25441 25594
rect 25441 25542 25453 25594
rect 25453 25542 25483 25594
rect 25507 25542 25517 25594
rect 25517 25542 25563 25594
rect 25267 25540 25323 25542
rect 25347 25540 25403 25542
rect 25427 25540 25483 25542
rect 25507 25540 25563 25542
rect 28354 25372 28356 25392
rect 28356 25372 28408 25392
rect 28408 25372 28410 25392
rect 28354 25336 28410 25372
rect 21794 25050 21850 25052
rect 21874 25050 21930 25052
rect 21954 25050 22010 25052
rect 22034 25050 22090 25052
rect 21794 24998 21840 25050
rect 21840 24998 21850 25050
rect 21874 24998 21904 25050
rect 21904 24998 21916 25050
rect 21916 24998 21930 25050
rect 21954 24998 21968 25050
rect 21968 24998 21980 25050
rect 21980 24998 22010 25050
rect 22034 24998 22044 25050
rect 22044 24998 22090 25050
rect 21794 24996 21850 24998
rect 21874 24996 21930 24998
rect 21954 24996 22010 24998
rect 22034 24996 22090 24998
rect 28740 25050 28796 25052
rect 28820 25050 28876 25052
rect 28900 25050 28956 25052
rect 28980 25050 29036 25052
rect 28740 24998 28786 25050
rect 28786 24998 28796 25050
rect 28820 24998 28850 25050
rect 28850 24998 28862 25050
rect 28862 24998 28876 25050
rect 28900 24998 28914 25050
rect 28914 24998 28926 25050
rect 28926 24998 28956 25050
rect 28980 24998 28990 25050
rect 28990 24998 29036 25050
rect 28740 24996 28796 24998
rect 28820 24996 28876 24998
rect 28900 24996 28956 24998
rect 28980 24996 29036 24998
rect 18321 24506 18377 24508
rect 18401 24506 18457 24508
rect 18481 24506 18537 24508
rect 18561 24506 18617 24508
rect 18321 24454 18367 24506
rect 18367 24454 18377 24506
rect 18401 24454 18431 24506
rect 18431 24454 18443 24506
rect 18443 24454 18457 24506
rect 18481 24454 18495 24506
rect 18495 24454 18507 24506
rect 18507 24454 18537 24506
rect 18561 24454 18571 24506
rect 18571 24454 18617 24506
rect 18321 24452 18377 24454
rect 18401 24452 18457 24454
rect 18481 24452 18537 24454
rect 18561 24452 18617 24454
rect 25267 24506 25323 24508
rect 25347 24506 25403 24508
rect 25427 24506 25483 24508
rect 25507 24506 25563 24508
rect 25267 24454 25313 24506
rect 25313 24454 25323 24506
rect 25347 24454 25377 24506
rect 25377 24454 25389 24506
rect 25389 24454 25403 24506
rect 25427 24454 25441 24506
rect 25441 24454 25453 24506
rect 25453 24454 25483 24506
rect 25507 24454 25517 24506
rect 25517 24454 25563 24506
rect 25267 24452 25323 24454
rect 25347 24452 25403 24454
rect 25427 24452 25483 24454
rect 25507 24452 25563 24454
rect 21794 23962 21850 23964
rect 21874 23962 21930 23964
rect 21954 23962 22010 23964
rect 22034 23962 22090 23964
rect 21794 23910 21840 23962
rect 21840 23910 21850 23962
rect 21874 23910 21904 23962
rect 21904 23910 21916 23962
rect 21916 23910 21930 23962
rect 21954 23910 21968 23962
rect 21968 23910 21980 23962
rect 21980 23910 22010 23962
rect 22034 23910 22044 23962
rect 22044 23910 22090 23962
rect 21794 23908 21850 23910
rect 21874 23908 21930 23910
rect 21954 23908 22010 23910
rect 22034 23908 22090 23910
rect 28740 23962 28796 23964
rect 28820 23962 28876 23964
rect 28900 23962 28956 23964
rect 28980 23962 29036 23964
rect 28740 23910 28786 23962
rect 28786 23910 28796 23962
rect 28820 23910 28850 23962
rect 28850 23910 28862 23962
rect 28862 23910 28876 23962
rect 28900 23910 28914 23962
rect 28914 23910 28926 23962
rect 28926 23910 28956 23962
rect 28980 23910 28990 23962
rect 28990 23910 29036 23962
rect 28740 23908 28796 23910
rect 28820 23908 28876 23910
rect 28900 23908 28956 23910
rect 28980 23908 29036 23910
rect 28354 23704 28410 23760
rect 18321 23418 18377 23420
rect 18401 23418 18457 23420
rect 18481 23418 18537 23420
rect 18561 23418 18617 23420
rect 18321 23366 18367 23418
rect 18367 23366 18377 23418
rect 18401 23366 18431 23418
rect 18431 23366 18443 23418
rect 18443 23366 18457 23418
rect 18481 23366 18495 23418
rect 18495 23366 18507 23418
rect 18507 23366 18537 23418
rect 18561 23366 18571 23418
rect 18571 23366 18617 23418
rect 18321 23364 18377 23366
rect 18401 23364 18457 23366
rect 18481 23364 18537 23366
rect 18561 23364 18617 23366
rect 25267 23418 25323 23420
rect 25347 23418 25403 23420
rect 25427 23418 25483 23420
rect 25507 23418 25563 23420
rect 25267 23366 25313 23418
rect 25313 23366 25323 23418
rect 25347 23366 25377 23418
rect 25377 23366 25389 23418
rect 25389 23366 25403 23418
rect 25427 23366 25441 23418
rect 25441 23366 25453 23418
rect 25453 23366 25483 23418
rect 25507 23366 25517 23418
rect 25517 23366 25563 23418
rect 25267 23364 25323 23366
rect 25347 23364 25403 23366
rect 25427 23364 25483 23366
rect 25507 23364 25563 23366
rect 28354 23060 28356 23080
rect 28356 23060 28408 23080
rect 28408 23060 28410 23080
rect 28354 23024 28410 23060
rect 21794 22874 21850 22876
rect 21874 22874 21930 22876
rect 21954 22874 22010 22876
rect 22034 22874 22090 22876
rect 21794 22822 21840 22874
rect 21840 22822 21850 22874
rect 21874 22822 21904 22874
rect 21904 22822 21916 22874
rect 21916 22822 21930 22874
rect 21954 22822 21968 22874
rect 21968 22822 21980 22874
rect 21980 22822 22010 22874
rect 22034 22822 22044 22874
rect 22044 22822 22090 22874
rect 21794 22820 21850 22822
rect 21874 22820 21930 22822
rect 21954 22820 22010 22822
rect 22034 22820 22090 22822
rect 28740 22874 28796 22876
rect 28820 22874 28876 22876
rect 28900 22874 28956 22876
rect 28980 22874 29036 22876
rect 28740 22822 28786 22874
rect 28786 22822 28796 22874
rect 28820 22822 28850 22874
rect 28850 22822 28862 22874
rect 28862 22822 28876 22874
rect 28900 22822 28914 22874
rect 28914 22822 28926 22874
rect 28926 22822 28956 22874
rect 28980 22822 28990 22874
rect 28990 22822 29036 22874
rect 28740 22820 28796 22822
rect 28820 22820 28876 22822
rect 28900 22820 28956 22822
rect 28980 22820 29036 22822
rect 18321 22330 18377 22332
rect 18401 22330 18457 22332
rect 18481 22330 18537 22332
rect 18561 22330 18617 22332
rect 18321 22278 18367 22330
rect 18367 22278 18377 22330
rect 18401 22278 18431 22330
rect 18431 22278 18443 22330
rect 18443 22278 18457 22330
rect 18481 22278 18495 22330
rect 18495 22278 18507 22330
rect 18507 22278 18537 22330
rect 18561 22278 18571 22330
rect 18571 22278 18617 22330
rect 18321 22276 18377 22278
rect 18401 22276 18457 22278
rect 18481 22276 18537 22278
rect 18561 22276 18617 22278
rect 25267 22330 25323 22332
rect 25347 22330 25403 22332
rect 25427 22330 25483 22332
rect 25507 22330 25563 22332
rect 25267 22278 25313 22330
rect 25313 22278 25323 22330
rect 25347 22278 25377 22330
rect 25377 22278 25389 22330
rect 25389 22278 25403 22330
rect 25427 22278 25441 22330
rect 25441 22278 25453 22330
rect 25453 22278 25483 22330
rect 25507 22278 25517 22330
rect 25517 22278 25563 22330
rect 25267 22276 25323 22278
rect 25347 22276 25403 22278
rect 25427 22276 25483 22278
rect 25507 22276 25563 22278
rect 28354 21972 28356 21992
rect 28356 21972 28408 21992
rect 28408 21972 28410 21992
rect 28354 21936 28410 21972
rect 21794 21786 21850 21788
rect 21874 21786 21930 21788
rect 21954 21786 22010 21788
rect 22034 21786 22090 21788
rect 21794 21734 21840 21786
rect 21840 21734 21850 21786
rect 21874 21734 21904 21786
rect 21904 21734 21916 21786
rect 21916 21734 21930 21786
rect 21954 21734 21968 21786
rect 21968 21734 21980 21786
rect 21980 21734 22010 21786
rect 22034 21734 22044 21786
rect 22044 21734 22090 21786
rect 21794 21732 21850 21734
rect 21874 21732 21930 21734
rect 21954 21732 22010 21734
rect 22034 21732 22090 21734
rect 28740 21786 28796 21788
rect 28820 21786 28876 21788
rect 28900 21786 28956 21788
rect 28980 21786 29036 21788
rect 28740 21734 28786 21786
rect 28786 21734 28796 21786
rect 28820 21734 28850 21786
rect 28850 21734 28862 21786
rect 28862 21734 28876 21786
rect 28900 21734 28914 21786
rect 28914 21734 28926 21786
rect 28926 21734 28956 21786
rect 28980 21734 28990 21786
rect 28990 21734 29036 21786
rect 28740 21732 28796 21734
rect 28820 21732 28876 21734
rect 28900 21732 28956 21734
rect 28980 21732 29036 21734
rect 18321 21242 18377 21244
rect 18401 21242 18457 21244
rect 18481 21242 18537 21244
rect 18561 21242 18617 21244
rect 18321 21190 18367 21242
rect 18367 21190 18377 21242
rect 18401 21190 18431 21242
rect 18431 21190 18443 21242
rect 18443 21190 18457 21242
rect 18481 21190 18495 21242
rect 18495 21190 18507 21242
rect 18507 21190 18537 21242
rect 18561 21190 18571 21242
rect 18571 21190 18617 21242
rect 18321 21188 18377 21190
rect 18401 21188 18457 21190
rect 18481 21188 18537 21190
rect 18561 21188 18617 21190
rect 25267 21242 25323 21244
rect 25347 21242 25403 21244
rect 25427 21242 25483 21244
rect 25507 21242 25563 21244
rect 25267 21190 25313 21242
rect 25313 21190 25323 21242
rect 25347 21190 25377 21242
rect 25377 21190 25389 21242
rect 25389 21190 25403 21242
rect 25427 21190 25441 21242
rect 25441 21190 25453 21242
rect 25453 21190 25483 21242
rect 25507 21190 25517 21242
rect 25517 21190 25563 21242
rect 25267 21188 25323 21190
rect 25347 21188 25403 21190
rect 25427 21188 25483 21190
rect 25507 21188 25563 21190
rect 28354 20984 28410 21040
rect 21794 20698 21850 20700
rect 21874 20698 21930 20700
rect 21954 20698 22010 20700
rect 22034 20698 22090 20700
rect 21794 20646 21840 20698
rect 21840 20646 21850 20698
rect 21874 20646 21904 20698
rect 21904 20646 21916 20698
rect 21916 20646 21930 20698
rect 21954 20646 21968 20698
rect 21968 20646 21980 20698
rect 21980 20646 22010 20698
rect 22034 20646 22044 20698
rect 22044 20646 22090 20698
rect 21794 20644 21850 20646
rect 21874 20644 21930 20646
rect 21954 20644 22010 20646
rect 22034 20644 22090 20646
rect 28740 20698 28796 20700
rect 28820 20698 28876 20700
rect 28900 20698 28956 20700
rect 28980 20698 29036 20700
rect 28740 20646 28786 20698
rect 28786 20646 28796 20698
rect 28820 20646 28850 20698
rect 28850 20646 28862 20698
rect 28862 20646 28876 20698
rect 28900 20646 28914 20698
rect 28914 20646 28926 20698
rect 28926 20646 28956 20698
rect 28980 20646 28990 20698
rect 28990 20646 29036 20698
rect 28740 20644 28796 20646
rect 28820 20644 28876 20646
rect 28900 20644 28956 20646
rect 28980 20644 29036 20646
rect 18321 20154 18377 20156
rect 18401 20154 18457 20156
rect 18481 20154 18537 20156
rect 18561 20154 18617 20156
rect 18321 20102 18367 20154
rect 18367 20102 18377 20154
rect 18401 20102 18431 20154
rect 18431 20102 18443 20154
rect 18443 20102 18457 20154
rect 18481 20102 18495 20154
rect 18495 20102 18507 20154
rect 18507 20102 18537 20154
rect 18561 20102 18571 20154
rect 18571 20102 18617 20154
rect 18321 20100 18377 20102
rect 18401 20100 18457 20102
rect 18481 20100 18537 20102
rect 18561 20100 18617 20102
rect 25267 20154 25323 20156
rect 25347 20154 25403 20156
rect 25427 20154 25483 20156
rect 25507 20154 25563 20156
rect 25267 20102 25313 20154
rect 25313 20102 25323 20154
rect 25347 20102 25377 20154
rect 25377 20102 25389 20154
rect 25389 20102 25403 20154
rect 25427 20102 25441 20154
rect 25441 20102 25453 20154
rect 25453 20102 25483 20154
rect 25507 20102 25517 20154
rect 25517 20102 25563 20154
rect 25267 20100 25323 20102
rect 25347 20100 25403 20102
rect 25427 20100 25483 20102
rect 25507 20100 25563 20102
rect 28354 19932 28356 19952
rect 28356 19932 28408 19952
rect 28408 19932 28410 19952
rect 28354 19896 28410 19932
rect 21794 19610 21850 19612
rect 21874 19610 21930 19612
rect 21954 19610 22010 19612
rect 22034 19610 22090 19612
rect 21794 19558 21840 19610
rect 21840 19558 21850 19610
rect 21874 19558 21904 19610
rect 21904 19558 21916 19610
rect 21916 19558 21930 19610
rect 21954 19558 21968 19610
rect 21968 19558 21980 19610
rect 21980 19558 22010 19610
rect 22034 19558 22044 19610
rect 22044 19558 22090 19610
rect 21794 19556 21850 19558
rect 21874 19556 21930 19558
rect 21954 19556 22010 19558
rect 22034 19556 22090 19558
rect 28740 19610 28796 19612
rect 28820 19610 28876 19612
rect 28900 19610 28956 19612
rect 28980 19610 29036 19612
rect 28740 19558 28786 19610
rect 28786 19558 28796 19610
rect 28820 19558 28850 19610
rect 28850 19558 28862 19610
rect 28862 19558 28876 19610
rect 28900 19558 28914 19610
rect 28914 19558 28926 19610
rect 28926 19558 28956 19610
rect 28980 19558 28990 19610
rect 28990 19558 29036 19610
rect 28740 19556 28796 19558
rect 28820 19556 28876 19558
rect 28900 19556 28956 19558
rect 28980 19556 29036 19558
rect 18321 19066 18377 19068
rect 18401 19066 18457 19068
rect 18481 19066 18537 19068
rect 18561 19066 18617 19068
rect 18321 19014 18367 19066
rect 18367 19014 18377 19066
rect 18401 19014 18431 19066
rect 18431 19014 18443 19066
rect 18443 19014 18457 19066
rect 18481 19014 18495 19066
rect 18495 19014 18507 19066
rect 18507 19014 18537 19066
rect 18561 19014 18571 19066
rect 18571 19014 18617 19066
rect 18321 19012 18377 19014
rect 18401 19012 18457 19014
rect 18481 19012 18537 19014
rect 18561 19012 18617 19014
rect 25267 19066 25323 19068
rect 25347 19066 25403 19068
rect 25427 19066 25483 19068
rect 25507 19066 25563 19068
rect 25267 19014 25313 19066
rect 25313 19014 25323 19066
rect 25347 19014 25377 19066
rect 25377 19014 25389 19066
rect 25389 19014 25403 19066
rect 25427 19014 25441 19066
rect 25441 19014 25453 19066
rect 25453 19014 25483 19066
rect 25507 19014 25517 19066
rect 25517 19014 25563 19066
rect 25267 19012 25323 19014
rect 25347 19012 25403 19014
rect 25427 19012 25483 19014
rect 25507 19012 25563 19014
rect 28354 18944 28410 19000
rect 21794 18522 21850 18524
rect 21874 18522 21930 18524
rect 21954 18522 22010 18524
rect 22034 18522 22090 18524
rect 21794 18470 21840 18522
rect 21840 18470 21850 18522
rect 21874 18470 21904 18522
rect 21904 18470 21916 18522
rect 21916 18470 21930 18522
rect 21954 18470 21968 18522
rect 21968 18470 21980 18522
rect 21980 18470 22010 18522
rect 22034 18470 22044 18522
rect 22044 18470 22090 18522
rect 21794 18468 21850 18470
rect 21874 18468 21930 18470
rect 21954 18468 22010 18470
rect 22034 18468 22090 18470
rect 28740 18522 28796 18524
rect 28820 18522 28876 18524
rect 28900 18522 28956 18524
rect 28980 18522 29036 18524
rect 28740 18470 28786 18522
rect 28786 18470 28796 18522
rect 28820 18470 28850 18522
rect 28850 18470 28862 18522
rect 28862 18470 28876 18522
rect 28900 18470 28914 18522
rect 28914 18470 28926 18522
rect 28926 18470 28956 18522
rect 28980 18470 28990 18522
rect 28990 18470 29036 18522
rect 28740 18468 28796 18470
rect 28820 18468 28876 18470
rect 28900 18468 28956 18470
rect 28980 18468 29036 18470
rect 18321 17978 18377 17980
rect 18401 17978 18457 17980
rect 18481 17978 18537 17980
rect 18561 17978 18617 17980
rect 18321 17926 18367 17978
rect 18367 17926 18377 17978
rect 18401 17926 18431 17978
rect 18431 17926 18443 17978
rect 18443 17926 18457 17978
rect 18481 17926 18495 17978
rect 18495 17926 18507 17978
rect 18507 17926 18537 17978
rect 18561 17926 18571 17978
rect 18571 17926 18617 17978
rect 18321 17924 18377 17926
rect 18401 17924 18457 17926
rect 18481 17924 18537 17926
rect 18561 17924 18617 17926
rect 25267 17978 25323 17980
rect 25347 17978 25403 17980
rect 25427 17978 25483 17980
rect 25507 17978 25563 17980
rect 25267 17926 25313 17978
rect 25313 17926 25323 17978
rect 25347 17926 25377 17978
rect 25377 17926 25389 17978
rect 25389 17926 25403 17978
rect 25427 17926 25441 17978
rect 25441 17926 25453 17978
rect 25453 17926 25483 17978
rect 25507 17926 25517 17978
rect 25517 17926 25563 17978
rect 25267 17924 25323 17926
rect 25347 17924 25403 17926
rect 25427 17924 25483 17926
rect 25507 17924 25563 17926
rect 28354 17620 28356 17640
rect 28356 17620 28408 17640
rect 28408 17620 28410 17640
rect 28354 17584 28410 17620
rect 21794 17434 21850 17436
rect 21874 17434 21930 17436
rect 21954 17434 22010 17436
rect 22034 17434 22090 17436
rect 21794 17382 21840 17434
rect 21840 17382 21850 17434
rect 21874 17382 21904 17434
rect 21904 17382 21916 17434
rect 21916 17382 21930 17434
rect 21954 17382 21968 17434
rect 21968 17382 21980 17434
rect 21980 17382 22010 17434
rect 22034 17382 22044 17434
rect 22044 17382 22090 17434
rect 21794 17380 21850 17382
rect 21874 17380 21930 17382
rect 21954 17380 22010 17382
rect 22034 17380 22090 17382
rect 28740 17434 28796 17436
rect 28820 17434 28876 17436
rect 28900 17434 28956 17436
rect 28980 17434 29036 17436
rect 28740 17382 28786 17434
rect 28786 17382 28796 17434
rect 28820 17382 28850 17434
rect 28850 17382 28862 17434
rect 28862 17382 28876 17434
rect 28900 17382 28914 17434
rect 28914 17382 28926 17434
rect 28926 17382 28956 17434
rect 28980 17382 28990 17434
rect 28990 17382 29036 17434
rect 28740 17380 28796 17382
rect 28820 17380 28876 17382
rect 28900 17380 28956 17382
rect 28980 17380 29036 17382
rect 28354 16940 28356 16960
rect 28356 16940 28408 16960
rect 28408 16940 28410 16960
rect 28354 16904 28410 16940
rect 18321 16890 18377 16892
rect 18401 16890 18457 16892
rect 18481 16890 18537 16892
rect 18561 16890 18617 16892
rect 18321 16838 18367 16890
rect 18367 16838 18377 16890
rect 18401 16838 18431 16890
rect 18431 16838 18443 16890
rect 18443 16838 18457 16890
rect 18481 16838 18495 16890
rect 18495 16838 18507 16890
rect 18507 16838 18537 16890
rect 18561 16838 18571 16890
rect 18571 16838 18617 16890
rect 18321 16836 18377 16838
rect 18401 16836 18457 16838
rect 18481 16836 18537 16838
rect 18561 16836 18617 16838
rect 25267 16890 25323 16892
rect 25347 16890 25403 16892
rect 25427 16890 25483 16892
rect 25507 16890 25563 16892
rect 25267 16838 25313 16890
rect 25313 16838 25323 16890
rect 25347 16838 25377 16890
rect 25377 16838 25389 16890
rect 25389 16838 25403 16890
rect 25427 16838 25441 16890
rect 25441 16838 25453 16890
rect 25453 16838 25483 16890
rect 25507 16838 25517 16890
rect 25517 16838 25563 16890
rect 25267 16836 25323 16838
rect 25347 16836 25403 16838
rect 25427 16836 25483 16838
rect 25507 16836 25563 16838
rect 21794 16346 21850 16348
rect 21874 16346 21930 16348
rect 21954 16346 22010 16348
rect 22034 16346 22090 16348
rect 21794 16294 21840 16346
rect 21840 16294 21850 16346
rect 21874 16294 21904 16346
rect 21904 16294 21916 16346
rect 21916 16294 21930 16346
rect 21954 16294 21968 16346
rect 21968 16294 21980 16346
rect 21980 16294 22010 16346
rect 22034 16294 22044 16346
rect 22044 16294 22090 16346
rect 21794 16292 21850 16294
rect 21874 16292 21930 16294
rect 21954 16292 22010 16294
rect 22034 16292 22090 16294
rect 28740 16346 28796 16348
rect 28820 16346 28876 16348
rect 28900 16346 28956 16348
rect 28980 16346 29036 16348
rect 28740 16294 28786 16346
rect 28786 16294 28796 16346
rect 28820 16294 28850 16346
rect 28850 16294 28862 16346
rect 28862 16294 28876 16346
rect 28900 16294 28914 16346
rect 28914 16294 28926 16346
rect 28926 16294 28956 16346
rect 28980 16294 28990 16346
rect 28990 16294 29036 16346
rect 28740 16292 28796 16294
rect 28820 16292 28876 16294
rect 28900 16292 28956 16294
rect 28980 16292 29036 16294
rect 18321 15802 18377 15804
rect 18401 15802 18457 15804
rect 18481 15802 18537 15804
rect 18561 15802 18617 15804
rect 18321 15750 18367 15802
rect 18367 15750 18377 15802
rect 18401 15750 18431 15802
rect 18431 15750 18443 15802
rect 18443 15750 18457 15802
rect 18481 15750 18495 15802
rect 18495 15750 18507 15802
rect 18507 15750 18537 15802
rect 18561 15750 18571 15802
rect 18571 15750 18617 15802
rect 18321 15748 18377 15750
rect 18401 15748 18457 15750
rect 18481 15748 18537 15750
rect 18561 15748 18617 15750
rect 25267 15802 25323 15804
rect 25347 15802 25403 15804
rect 25427 15802 25483 15804
rect 25507 15802 25563 15804
rect 25267 15750 25313 15802
rect 25313 15750 25323 15802
rect 25347 15750 25377 15802
rect 25377 15750 25389 15802
rect 25389 15750 25403 15802
rect 25427 15750 25441 15802
rect 25441 15750 25453 15802
rect 25453 15750 25483 15802
rect 25507 15750 25517 15802
rect 25517 15750 25563 15802
rect 25267 15748 25323 15750
rect 25347 15748 25403 15750
rect 25427 15748 25483 15750
rect 25507 15748 25563 15750
rect 28354 15544 28410 15600
rect 21794 15258 21850 15260
rect 21874 15258 21930 15260
rect 21954 15258 22010 15260
rect 22034 15258 22090 15260
rect 21794 15206 21840 15258
rect 21840 15206 21850 15258
rect 21874 15206 21904 15258
rect 21904 15206 21916 15258
rect 21916 15206 21930 15258
rect 21954 15206 21968 15258
rect 21968 15206 21980 15258
rect 21980 15206 22010 15258
rect 22034 15206 22044 15258
rect 22044 15206 22090 15258
rect 21794 15204 21850 15206
rect 21874 15204 21930 15206
rect 21954 15204 22010 15206
rect 22034 15204 22090 15206
rect 28740 15258 28796 15260
rect 28820 15258 28876 15260
rect 28900 15258 28956 15260
rect 28980 15258 29036 15260
rect 28740 15206 28786 15258
rect 28786 15206 28796 15258
rect 28820 15206 28850 15258
rect 28850 15206 28862 15258
rect 28862 15206 28876 15258
rect 28900 15206 28914 15258
rect 28914 15206 28926 15258
rect 28926 15206 28956 15258
rect 28980 15206 28990 15258
rect 28990 15206 29036 15258
rect 28740 15204 28796 15206
rect 28820 15204 28876 15206
rect 28900 15204 28956 15206
rect 28980 15204 29036 15206
rect 28354 14884 28410 14920
rect 28354 14864 28356 14884
rect 28356 14864 28408 14884
rect 28408 14864 28410 14884
rect 18321 14714 18377 14716
rect 18401 14714 18457 14716
rect 18481 14714 18537 14716
rect 18561 14714 18617 14716
rect 18321 14662 18367 14714
rect 18367 14662 18377 14714
rect 18401 14662 18431 14714
rect 18431 14662 18443 14714
rect 18443 14662 18457 14714
rect 18481 14662 18495 14714
rect 18495 14662 18507 14714
rect 18507 14662 18537 14714
rect 18561 14662 18571 14714
rect 18571 14662 18617 14714
rect 18321 14660 18377 14662
rect 18401 14660 18457 14662
rect 18481 14660 18537 14662
rect 18561 14660 18617 14662
rect 25267 14714 25323 14716
rect 25347 14714 25403 14716
rect 25427 14714 25483 14716
rect 25507 14714 25563 14716
rect 25267 14662 25313 14714
rect 25313 14662 25323 14714
rect 25347 14662 25377 14714
rect 25377 14662 25389 14714
rect 25389 14662 25403 14714
rect 25427 14662 25441 14714
rect 25441 14662 25453 14714
rect 25453 14662 25483 14714
rect 25507 14662 25517 14714
rect 25517 14662 25563 14714
rect 25267 14660 25323 14662
rect 25347 14660 25403 14662
rect 25427 14660 25483 14662
rect 25507 14660 25563 14662
rect 21794 14170 21850 14172
rect 21874 14170 21930 14172
rect 21954 14170 22010 14172
rect 22034 14170 22090 14172
rect 21794 14118 21840 14170
rect 21840 14118 21850 14170
rect 21874 14118 21904 14170
rect 21904 14118 21916 14170
rect 21916 14118 21930 14170
rect 21954 14118 21968 14170
rect 21968 14118 21980 14170
rect 21980 14118 22010 14170
rect 22034 14118 22044 14170
rect 22044 14118 22090 14170
rect 21794 14116 21850 14118
rect 21874 14116 21930 14118
rect 21954 14116 22010 14118
rect 22034 14116 22090 14118
rect 28740 14170 28796 14172
rect 28820 14170 28876 14172
rect 28900 14170 28956 14172
rect 28980 14170 29036 14172
rect 28740 14118 28786 14170
rect 28786 14118 28796 14170
rect 28820 14118 28850 14170
rect 28850 14118 28862 14170
rect 28862 14118 28876 14170
rect 28900 14118 28914 14170
rect 28914 14118 28926 14170
rect 28926 14118 28956 14170
rect 28980 14118 28990 14170
rect 28990 14118 29036 14170
rect 28740 14116 28796 14118
rect 28820 14116 28876 14118
rect 28900 14116 28956 14118
rect 28980 14116 29036 14118
rect 18321 13626 18377 13628
rect 18401 13626 18457 13628
rect 18481 13626 18537 13628
rect 18561 13626 18617 13628
rect 18321 13574 18367 13626
rect 18367 13574 18377 13626
rect 18401 13574 18431 13626
rect 18431 13574 18443 13626
rect 18443 13574 18457 13626
rect 18481 13574 18495 13626
rect 18495 13574 18507 13626
rect 18507 13574 18537 13626
rect 18561 13574 18571 13626
rect 18571 13574 18617 13626
rect 18321 13572 18377 13574
rect 18401 13572 18457 13574
rect 18481 13572 18537 13574
rect 18561 13572 18617 13574
rect 25267 13626 25323 13628
rect 25347 13626 25403 13628
rect 25427 13626 25483 13628
rect 25507 13626 25563 13628
rect 25267 13574 25313 13626
rect 25313 13574 25323 13626
rect 25347 13574 25377 13626
rect 25377 13574 25389 13626
rect 25389 13574 25403 13626
rect 25427 13574 25441 13626
rect 25441 13574 25453 13626
rect 25453 13574 25483 13626
rect 25507 13574 25517 13626
rect 25517 13574 25563 13626
rect 25267 13572 25323 13574
rect 25347 13572 25403 13574
rect 25427 13572 25483 13574
rect 25507 13572 25563 13574
rect 28354 13504 28410 13560
rect 21794 13082 21850 13084
rect 21874 13082 21930 13084
rect 21954 13082 22010 13084
rect 22034 13082 22090 13084
rect 21794 13030 21840 13082
rect 21840 13030 21850 13082
rect 21874 13030 21904 13082
rect 21904 13030 21916 13082
rect 21916 13030 21930 13082
rect 21954 13030 21968 13082
rect 21968 13030 21980 13082
rect 21980 13030 22010 13082
rect 22034 13030 22044 13082
rect 22044 13030 22090 13082
rect 21794 13028 21850 13030
rect 21874 13028 21930 13030
rect 21954 13028 22010 13030
rect 22034 13028 22090 13030
rect 28740 13082 28796 13084
rect 28820 13082 28876 13084
rect 28900 13082 28956 13084
rect 28980 13082 29036 13084
rect 28740 13030 28786 13082
rect 28786 13030 28796 13082
rect 28820 13030 28850 13082
rect 28850 13030 28862 13082
rect 28862 13030 28876 13082
rect 28900 13030 28914 13082
rect 28914 13030 28926 13082
rect 28926 13030 28956 13082
rect 28980 13030 28990 13082
rect 28990 13030 29036 13082
rect 28740 13028 28796 13030
rect 28820 13028 28876 13030
rect 28900 13028 28956 13030
rect 28980 13028 29036 13030
rect 28354 12824 28410 12880
rect 18321 12538 18377 12540
rect 18401 12538 18457 12540
rect 18481 12538 18537 12540
rect 18561 12538 18617 12540
rect 18321 12486 18367 12538
rect 18367 12486 18377 12538
rect 18401 12486 18431 12538
rect 18431 12486 18443 12538
rect 18443 12486 18457 12538
rect 18481 12486 18495 12538
rect 18495 12486 18507 12538
rect 18507 12486 18537 12538
rect 18561 12486 18571 12538
rect 18571 12486 18617 12538
rect 18321 12484 18377 12486
rect 18401 12484 18457 12486
rect 18481 12484 18537 12486
rect 18561 12484 18617 12486
rect 25267 12538 25323 12540
rect 25347 12538 25403 12540
rect 25427 12538 25483 12540
rect 25507 12538 25563 12540
rect 25267 12486 25313 12538
rect 25313 12486 25323 12538
rect 25347 12486 25377 12538
rect 25377 12486 25389 12538
rect 25389 12486 25403 12538
rect 25427 12486 25441 12538
rect 25441 12486 25453 12538
rect 25453 12486 25483 12538
rect 25507 12486 25517 12538
rect 25517 12486 25563 12538
rect 25267 12484 25323 12486
rect 25347 12484 25403 12486
rect 25427 12484 25483 12486
rect 25507 12484 25563 12486
rect 21794 11994 21850 11996
rect 21874 11994 21930 11996
rect 21954 11994 22010 11996
rect 22034 11994 22090 11996
rect 21794 11942 21840 11994
rect 21840 11942 21850 11994
rect 21874 11942 21904 11994
rect 21904 11942 21916 11994
rect 21916 11942 21930 11994
rect 21954 11942 21968 11994
rect 21968 11942 21980 11994
rect 21980 11942 22010 11994
rect 22034 11942 22044 11994
rect 22044 11942 22090 11994
rect 21794 11940 21850 11942
rect 21874 11940 21930 11942
rect 21954 11940 22010 11942
rect 22034 11940 22090 11942
rect 28740 11994 28796 11996
rect 28820 11994 28876 11996
rect 28900 11994 28956 11996
rect 28980 11994 29036 11996
rect 28740 11942 28786 11994
rect 28786 11942 28796 11994
rect 28820 11942 28850 11994
rect 28850 11942 28862 11994
rect 28862 11942 28876 11994
rect 28900 11942 28914 11994
rect 28914 11942 28926 11994
rect 28926 11942 28956 11994
rect 28980 11942 28990 11994
rect 28990 11942 29036 11994
rect 28740 11940 28796 11942
rect 28820 11940 28876 11942
rect 28900 11940 28956 11942
rect 28980 11940 29036 11942
rect 28354 11500 28356 11520
rect 28356 11500 28408 11520
rect 28408 11500 28410 11520
rect 28354 11464 28410 11500
rect 18321 11450 18377 11452
rect 18401 11450 18457 11452
rect 18481 11450 18537 11452
rect 18561 11450 18617 11452
rect 18321 11398 18367 11450
rect 18367 11398 18377 11450
rect 18401 11398 18431 11450
rect 18431 11398 18443 11450
rect 18443 11398 18457 11450
rect 18481 11398 18495 11450
rect 18495 11398 18507 11450
rect 18507 11398 18537 11450
rect 18561 11398 18571 11450
rect 18571 11398 18617 11450
rect 18321 11396 18377 11398
rect 18401 11396 18457 11398
rect 18481 11396 18537 11398
rect 18561 11396 18617 11398
rect 25267 11450 25323 11452
rect 25347 11450 25403 11452
rect 25427 11450 25483 11452
rect 25507 11450 25563 11452
rect 25267 11398 25313 11450
rect 25313 11398 25323 11450
rect 25347 11398 25377 11450
rect 25377 11398 25389 11450
rect 25389 11398 25403 11450
rect 25427 11398 25441 11450
rect 25441 11398 25453 11450
rect 25453 11398 25483 11450
rect 25507 11398 25517 11450
rect 25517 11398 25563 11450
rect 25267 11396 25323 11398
rect 25347 11396 25403 11398
rect 25427 11396 25483 11398
rect 25507 11396 25563 11398
rect 28354 11092 28356 11112
rect 28356 11092 28408 11112
rect 28408 11092 28410 11112
rect 28354 11056 28410 11092
rect 21794 10906 21850 10908
rect 21874 10906 21930 10908
rect 21954 10906 22010 10908
rect 22034 10906 22090 10908
rect 21794 10854 21840 10906
rect 21840 10854 21850 10906
rect 21874 10854 21904 10906
rect 21904 10854 21916 10906
rect 21916 10854 21930 10906
rect 21954 10854 21968 10906
rect 21968 10854 21980 10906
rect 21980 10854 22010 10906
rect 22034 10854 22044 10906
rect 22044 10854 22090 10906
rect 21794 10852 21850 10854
rect 21874 10852 21930 10854
rect 21954 10852 22010 10854
rect 22034 10852 22090 10854
rect 28740 10906 28796 10908
rect 28820 10906 28876 10908
rect 28900 10906 28956 10908
rect 28980 10906 29036 10908
rect 28740 10854 28786 10906
rect 28786 10854 28796 10906
rect 28820 10854 28850 10906
rect 28850 10854 28862 10906
rect 28862 10854 28876 10906
rect 28900 10854 28914 10906
rect 28914 10854 28926 10906
rect 28926 10854 28956 10906
rect 28980 10854 28990 10906
rect 28990 10854 29036 10906
rect 28740 10852 28796 10854
rect 28820 10852 28876 10854
rect 28900 10852 28956 10854
rect 28980 10852 29036 10854
rect 18321 10362 18377 10364
rect 18401 10362 18457 10364
rect 18481 10362 18537 10364
rect 18561 10362 18617 10364
rect 18321 10310 18367 10362
rect 18367 10310 18377 10362
rect 18401 10310 18431 10362
rect 18431 10310 18443 10362
rect 18443 10310 18457 10362
rect 18481 10310 18495 10362
rect 18495 10310 18507 10362
rect 18507 10310 18537 10362
rect 18561 10310 18571 10362
rect 18571 10310 18617 10362
rect 18321 10308 18377 10310
rect 18401 10308 18457 10310
rect 18481 10308 18537 10310
rect 18561 10308 18617 10310
rect 25267 10362 25323 10364
rect 25347 10362 25403 10364
rect 25427 10362 25483 10364
rect 25507 10362 25563 10364
rect 25267 10310 25313 10362
rect 25313 10310 25323 10362
rect 25347 10310 25377 10362
rect 25377 10310 25389 10362
rect 25389 10310 25403 10362
rect 25427 10310 25441 10362
rect 25441 10310 25453 10362
rect 25453 10310 25483 10362
rect 25507 10310 25517 10362
rect 25517 10310 25563 10362
rect 25267 10308 25323 10310
rect 25347 10308 25403 10310
rect 25427 10308 25483 10310
rect 25507 10308 25563 10310
rect 21794 9818 21850 9820
rect 21874 9818 21930 9820
rect 21954 9818 22010 9820
rect 22034 9818 22090 9820
rect 21794 9766 21840 9818
rect 21840 9766 21850 9818
rect 21874 9766 21904 9818
rect 21904 9766 21916 9818
rect 21916 9766 21930 9818
rect 21954 9766 21968 9818
rect 21968 9766 21980 9818
rect 21980 9766 22010 9818
rect 22034 9766 22044 9818
rect 22044 9766 22090 9818
rect 21794 9764 21850 9766
rect 21874 9764 21930 9766
rect 21954 9764 22010 9766
rect 22034 9764 22090 9766
rect 28740 9818 28796 9820
rect 28820 9818 28876 9820
rect 28900 9818 28956 9820
rect 28980 9818 29036 9820
rect 28740 9766 28786 9818
rect 28786 9766 28796 9818
rect 28820 9766 28850 9818
rect 28850 9766 28862 9818
rect 28862 9766 28876 9818
rect 28900 9766 28914 9818
rect 28914 9766 28926 9818
rect 28926 9766 28956 9818
rect 28980 9766 28990 9818
rect 28990 9766 29036 9818
rect 28740 9764 28796 9766
rect 28820 9764 28876 9766
rect 28900 9764 28956 9766
rect 28980 9764 29036 9766
rect 28354 9444 28410 9480
rect 28354 9424 28356 9444
rect 28356 9424 28408 9444
rect 28408 9424 28410 9444
rect 18321 9274 18377 9276
rect 18401 9274 18457 9276
rect 18481 9274 18537 9276
rect 18561 9274 18617 9276
rect 18321 9222 18367 9274
rect 18367 9222 18377 9274
rect 18401 9222 18431 9274
rect 18431 9222 18443 9274
rect 18443 9222 18457 9274
rect 18481 9222 18495 9274
rect 18495 9222 18507 9274
rect 18507 9222 18537 9274
rect 18561 9222 18571 9274
rect 18571 9222 18617 9274
rect 18321 9220 18377 9222
rect 18401 9220 18457 9222
rect 18481 9220 18537 9222
rect 18561 9220 18617 9222
rect 25267 9274 25323 9276
rect 25347 9274 25403 9276
rect 25427 9274 25483 9276
rect 25507 9274 25563 9276
rect 25267 9222 25313 9274
rect 25313 9222 25323 9274
rect 25347 9222 25377 9274
rect 25377 9222 25389 9274
rect 25389 9222 25403 9274
rect 25427 9222 25441 9274
rect 25441 9222 25453 9274
rect 25453 9222 25483 9274
rect 25507 9222 25517 9274
rect 25517 9222 25563 9274
rect 25267 9220 25323 9222
rect 25347 9220 25403 9222
rect 25427 9220 25483 9222
rect 25507 9220 25563 9222
rect 28354 9052 28356 9072
rect 28356 9052 28408 9072
rect 28408 9052 28410 9072
rect 28354 9016 28410 9052
rect 21794 8730 21850 8732
rect 21874 8730 21930 8732
rect 21954 8730 22010 8732
rect 22034 8730 22090 8732
rect 21794 8678 21840 8730
rect 21840 8678 21850 8730
rect 21874 8678 21904 8730
rect 21904 8678 21916 8730
rect 21916 8678 21930 8730
rect 21954 8678 21968 8730
rect 21968 8678 21980 8730
rect 21980 8678 22010 8730
rect 22034 8678 22044 8730
rect 22044 8678 22090 8730
rect 21794 8676 21850 8678
rect 21874 8676 21930 8678
rect 21954 8676 22010 8678
rect 22034 8676 22090 8678
rect 28740 8730 28796 8732
rect 28820 8730 28876 8732
rect 28900 8730 28956 8732
rect 28980 8730 29036 8732
rect 28740 8678 28786 8730
rect 28786 8678 28796 8730
rect 28820 8678 28850 8730
rect 28850 8678 28862 8730
rect 28862 8678 28876 8730
rect 28900 8678 28914 8730
rect 28914 8678 28926 8730
rect 28926 8678 28956 8730
rect 28980 8678 28990 8730
rect 28990 8678 29036 8730
rect 28740 8676 28796 8678
rect 28820 8676 28876 8678
rect 28900 8676 28956 8678
rect 28980 8676 29036 8678
rect 18321 8186 18377 8188
rect 18401 8186 18457 8188
rect 18481 8186 18537 8188
rect 18561 8186 18617 8188
rect 18321 8134 18367 8186
rect 18367 8134 18377 8186
rect 18401 8134 18431 8186
rect 18431 8134 18443 8186
rect 18443 8134 18457 8186
rect 18481 8134 18495 8186
rect 18495 8134 18507 8186
rect 18507 8134 18537 8186
rect 18561 8134 18571 8186
rect 18571 8134 18617 8186
rect 18321 8132 18377 8134
rect 18401 8132 18457 8134
rect 18481 8132 18537 8134
rect 18561 8132 18617 8134
rect 25267 8186 25323 8188
rect 25347 8186 25403 8188
rect 25427 8186 25483 8188
rect 25507 8186 25563 8188
rect 25267 8134 25313 8186
rect 25313 8134 25323 8186
rect 25347 8134 25377 8186
rect 25377 8134 25389 8186
rect 25389 8134 25403 8186
rect 25427 8134 25441 8186
rect 25441 8134 25453 8186
rect 25453 8134 25483 8186
rect 25507 8134 25517 8186
rect 25517 8134 25563 8186
rect 25267 8132 25323 8134
rect 25347 8132 25403 8134
rect 25427 8132 25483 8134
rect 25507 8132 25563 8134
rect 21794 7642 21850 7644
rect 21874 7642 21930 7644
rect 21954 7642 22010 7644
rect 22034 7642 22090 7644
rect 21794 7590 21840 7642
rect 21840 7590 21850 7642
rect 21874 7590 21904 7642
rect 21904 7590 21916 7642
rect 21916 7590 21930 7642
rect 21954 7590 21968 7642
rect 21968 7590 21980 7642
rect 21980 7590 22010 7642
rect 22034 7590 22044 7642
rect 22044 7590 22090 7642
rect 21794 7588 21850 7590
rect 21874 7588 21930 7590
rect 21954 7588 22010 7590
rect 22034 7588 22090 7590
rect 28740 7642 28796 7644
rect 28820 7642 28876 7644
rect 28900 7642 28956 7644
rect 28980 7642 29036 7644
rect 28740 7590 28786 7642
rect 28786 7590 28796 7642
rect 28820 7590 28850 7642
rect 28850 7590 28862 7642
rect 28862 7590 28876 7642
rect 28900 7590 28914 7642
rect 28914 7590 28926 7642
rect 28926 7590 28956 7642
rect 28980 7590 28990 7642
rect 28990 7590 29036 7642
rect 28740 7588 28796 7590
rect 28820 7588 28876 7590
rect 28900 7588 28956 7590
rect 28980 7588 29036 7590
rect 28354 7384 28410 7440
rect 18321 7098 18377 7100
rect 18401 7098 18457 7100
rect 18481 7098 18537 7100
rect 18561 7098 18617 7100
rect 18321 7046 18367 7098
rect 18367 7046 18377 7098
rect 18401 7046 18431 7098
rect 18431 7046 18443 7098
rect 18443 7046 18457 7098
rect 18481 7046 18495 7098
rect 18495 7046 18507 7098
rect 18507 7046 18537 7098
rect 18561 7046 18571 7098
rect 18571 7046 18617 7098
rect 18321 7044 18377 7046
rect 18401 7044 18457 7046
rect 18481 7044 18537 7046
rect 18561 7044 18617 7046
rect 25267 7098 25323 7100
rect 25347 7098 25403 7100
rect 25427 7098 25483 7100
rect 25507 7098 25563 7100
rect 25267 7046 25313 7098
rect 25313 7046 25323 7098
rect 25347 7046 25377 7098
rect 25377 7046 25389 7098
rect 25389 7046 25403 7098
rect 25427 7046 25441 7098
rect 25441 7046 25453 7098
rect 25453 7046 25483 7098
rect 25507 7046 25517 7098
rect 25517 7046 25563 7098
rect 25267 7044 25323 7046
rect 25347 7044 25403 7046
rect 25427 7044 25483 7046
rect 25507 7044 25563 7046
rect 28354 6740 28356 6760
rect 28356 6740 28408 6760
rect 28408 6740 28410 6760
rect 28354 6704 28410 6740
rect 21794 6554 21850 6556
rect 21874 6554 21930 6556
rect 21954 6554 22010 6556
rect 22034 6554 22090 6556
rect 21794 6502 21840 6554
rect 21840 6502 21850 6554
rect 21874 6502 21904 6554
rect 21904 6502 21916 6554
rect 21916 6502 21930 6554
rect 21954 6502 21968 6554
rect 21968 6502 21980 6554
rect 21980 6502 22010 6554
rect 22034 6502 22044 6554
rect 22044 6502 22090 6554
rect 21794 6500 21850 6502
rect 21874 6500 21930 6502
rect 21954 6500 22010 6502
rect 22034 6500 22090 6502
rect 28740 6554 28796 6556
rect 28820 6554 28876 6556
rect 28900 6554 28956 6556
rect 28980 6554 29036 6556
rect 28740 6502 28786 6554
rect 28786 6502 28796 6554
rect 28820 6502 28850 6554
rect 28850 6502 28862 6554
rect 28862 6502 28876 6554
rect 28900 6502 28914 6554
rect 28914 6502 28926 6554
rect 28926 6502 28956 6554
rect 28980 6502 28990 6554
rect 28990 6502 29036 6554
rect 28740 6500 28796 6502
rect 28820 6500 28876 6502
rect 28900 6500 28956 6502
rect 28980 6500 29036 6502
rect 18321 6010 18377 6012
rect 18401 6010 18457 6012
rect 18481 6010 18537 6012
rect 18561 6010 18617 6012
rect 18321 5958 18367 6010
rect 18367 5958 18377 6010
rect 18401 5958 18431 6010
rect 18431 5958 18443 6010
rect 18443 5958 18457 6010
rect 18481 5958 18495 6010
rect 18495 5958 18507 6010
rect 18507 5958 18537 6010
rect 18561 5958 18571 6010
rect 18571 5958 18617 6010
rect 18321 5956 18377 5958
rect 18401 5956 18457 5958
rect 18481 5956 18537 5958
rect 18561 5956 18617 5958
rect 25267 6010 25323 6012
rect 25347 6010 25403 6012
rect 25427 6010 25483 6012
rect 25507 6010 25563 6012
rect 25267 5958 25313 6010
rect 25313 5958 25323 6010
rect 25347 5958 25377 6010
rect 25377 5958 25389 6010
rect 25389 5958 25403 6010
rect 25427 5958 25441 6010
rect 25441 5958 25453 6010
rect 25453 5958 25483 6010
rect 25507 5958 25517 6010
rect 25517 5958 25563 6010
rect 25267 5956 25323 5958
rect 25347 5956 25403 5958
rect 25427 5956 25483 5958
rect 25507 5956 25563 5958
rect 28354 5652 28356 5672
rect 28356 5652 28408 5672
rect 28408 5652 28410 5672
rect 28354 5616 28410 5652
rect 21794 5466 21850 5468
rect 21874 5466 21930 5468
rect 21954 5466 22010 5468
rect 22034 5466 22090 5468
rect 21794 5414 21840 5466
rect 21840 5414 21850 5466
rect 21874 5414 21904 5466
rect 21904 5414 21916 5466
rect 21916 5414 21930 5466
rect 21954 5414 21968 5466
rect 21968 5414 21980 5466
rect 21980 5414 22010 5466
rect 22034 5414 22044 5466
rect 22044 5414 22090 5466
rect 21794 5412 21850 5414
rect 21874 5412 21930 5414
rect 21954 5412 22010 5414
rect 22034 5412 22090 5414
rect 28740 5466 28796 5468
rect 28820 5466 28876 5468
rect 28900 5466 28956 5468
rect 28980 5466 29036 5468
rect 28740 5414 28786 5466
rect 28786 5414 28796 5466
rect 28820 5414 28850 5466
rect 28850 5414 28862 5466
rect 28862 5414 28876 5466
rect 28900 5414 28914 5466
rect 28914 5414 28926 5466
rect 28926 5414 28956 5466
rect 28980 5414 28990 5466
rect 28990 5414 29036 5466
rect 28740 5412 28796 5414
rect 28820 5412 28876 5414
rect 28900 5412 28956 5414
rect 28980 5412 29036 5414
rect 18321 4922 18377 4924
rect 18401 4922 18457 4924
rect 18481 4922 18537 4924
rect 18561 4922 18617 4924
rect 18321 4870 18367 4922
rect 18367 4870 18377 4922
rect 18401 4870 18431 4922
rect 18431 4870 18443 4922
rect 18443 4870 18457 4922
rect 18481 4870 18495 4922
rect 18495 4870 18507 4922
rect 18507 4870 18537 4922
rect 18561 4870 18571 4922
rect 18571 4870 18617 4922
rect 18321 4868 18377 4870
rect 18401 4868 18457 4870
rect 18481 4868 18537 4870
rect 18561 4868 18617 4870
rect 25267 4922 25323 4924
rect 25347 4922 25403 4924
rect 25427 4922 25483 4924
rect 25507 4922 25563 4924
rect 25267 4870 25313 4922
rect 25313 4870 25323 4922
rect 25347 4870 25377 4922
rect 25377 4870 25389 4922
rect 25389 4870 25403 4922
rect 25427 4870 25441 4922
rect 25441 4870 25453 4922
rect 25453 4870 25483 4922
rect 25507 4870 25517 4922
rect 25517 4870 25563 4922
rect 25267 4868 25323 4870
rect 25347 4868 25403 4870
rect 25427 4868 25483 4870
rect 25507 4868 25563 4870
rect 28354 4664 28410 4720
rect 21794 4378 21850 4380
rect 21874 4378 21930 4380
rect 21954 4378 22010 4380
rect 22034 4378 22090 4380
rect 21794 4326 21840 4378
rect 21840 4326 21850 4378
rect 21874 4326 21904 4378
rect 21904 4326 21916 4378
rect 21916 4326 21930 4378
rect 21954 4326 21968 4378
rect 21968 4326 21980 4378
rect 21980 4326 22010 4378
rect 22034 4326 22044 4378
rect 22044 4326 22090 4378
rect 21794 4324 21850 4326
rect 21874 4324 21930 4326
rect 21954 4324 22010 4326
rect 22034 4324 22090 4326
rect 28740 4378 28796 4380
rect 28820 4378 28876 4380
rect 28900 4378 28956 4380
rect 28980 4378 29036 4380
rect 28740 4326 28786 4378
rect 28786 4326 28796 4378
rect 28820 4326 28850 4378
rect 28850 4326 28862 4378
rect 28862 4326 28876 4378
rect 28900 4326 28914 4378
rect 28914 4326 28926 4378
rect 28926 4326 28956 4378
rect 28980 4326 28990 4378
rect 28990 4326 29036 4378
rect 28740 4324 28796 4326
rect 28820 4324 28876 4326
rect 28900 4324 28956 4326
rect 28980 4324 29036 4326
rect 28354 4020 28356 4040
rect 28356 4020 28408 4040
rect 28408 4020 28410 4040
rect 28354 3984 28410 4020
rect 4429 3834 4485 3836
rect 4509 3834 4565 3836
rect 4589 3834 4645 3836
rect 4669 3834 4725 3836
rect 4429 3782 4475 3834
rect 4475 3782 4485 3834
rect 4509 3782 4539 3834
rect 4539 3782 4551 3834
rect 4551 3782 4565 3834
rect 4589 3782 4603 3834
rect 4603 3782 4615 3834
rect 4615 3782 4645 3834
rect 4669 3782 4679 3834
rect 4679 3782 4725 3834
rect 4429 3780 4485 3782
rect 4509 3780 4565 3782
rect 4589 3780 4645 3782
rect 4669 3780 4725 3782
rect 11375 3834 11431 3836
rect 11455 3834 11511 3836
rect 11535 3834 11591 3836
rect 11615 3834 11671 3836
rect 11375 3782 11421 3834
rect 11421 3782 11431 3834
rect 11455 3782 11485 3834
rect 11485 3782 11497 3834
rect 11497 3782 11511 3834
rect 11535 3782 11549 3834
rect 11549 3782 11561 3834
rect 11561 3782 11591 3834
rect 11615 3782 11625 3834
rect 11625 3782 11671 3834
rect 11375 3780 11431 3782
rect 11455 3780 11511 3782
rect 11535 3780 11591 3782
rect 11615 3780 11671 3782
rect 18321 3834 18377 3836
rect 18401 3834 18457 3836
rect 18481 3834 18537 3836
rect 18561 3834 18617 3836
rect 18321 3782 18367 3834
rect 18367 3782 18377 3834
rect 18401 3782 18431 3834
rect 18431 3782 18443 3834
rect 18443 3782 18457 3834
rect 18481 3782 18495 3834
rect 18495 3782 18507 3834
rect 18507 3782 18537 3834
rect 18561 3782 18571 3834
rect 18571 3782 18617 3834
rect 18321 3780 18377 3782
rect 18401 3780 18457 3782
rect 18481 3780 18537 3782
rect 18561 3780 18617 3782
rect 25267 3834 25323 3836
rect 25347 3834 25403 3836
rect 25427 3834 25483 3836
rect 25507 3834 25563 3836
rect 25267 3782 25313 3834
rect 25313 3782 25323 3834
rect 25347 3782 25377 3834
rect 25377 3782 25389 3834
rect 25389 3782 25403 3834
rect 25427 3782 25441 3834
rect 25441 3782 25453 3834
rect 25453 3782 25483 3834
rect 25507 3782 25517 3834
rect 25517 3782 25563 3834
rect 25267 3780 25323 3782
rect 25347 3780 25403 3782
rect 25427 3780 25483 3782
rect 25507 3780 25563 3782
rect 1582 3712 1638 3768
rect 28354 3612 28356 3632
rect 28356 3612 28408 3632
rect 28408 3612 28410 3632
rect 28354 3576 28410 3612
rect 7902 3290 7958 3292
rect 7982 3290 8038 3292
rect 8062 3290 8118 3292
rect 8142 3290 8198 3292
rect 7902 3238 7948 3290
rect 7948 3238 7958 3290
rect 7982 3238 8012 3290
rect 8012 3238 8024 3290
rect 8024 3238 8038 3290
rect 8062 3238 8076 3290
rect 8076 3238 8088 3290
rect 8088 3238 8118 3290
rect 8142 3238 8152 3290
rect 8152 3238 8198 3290
rect 7902 3236 7958 3238
rect 7982 3236 8038 3238
rect 8062 3236 8118 3238
rect 8142 3236 8198 3238
rect 14848 3290 14904 3292
rect 14928 3290 14984 3292
rect 15008 3290 15064 3292
rect 15088 3290 15144 3292
rect 14848 3238 14894 3290
rect 14894 3238 14904 3290
rect 14928 3238 14958 3290
rect 14958 3238 14970 3290
rect 14970 3238 14984 3290
rect 15008 3238 15022 3290
rect 15022 3238 15034 3290
rect 15034 3238 15064 3290
rect 15088 3238 15098 3290
rect 15098 3238 15144 3290
rect 14848 3236 14904 3238
rect 14928 3236 14984 3238
rect 15008 3236 15064 3238
rect 15088 3236 15144 3238
rect 21794 3290 21850 3292
rect 21874 3290 21930 3292
rect 21954 3290 22010 3292
rect 22034 3290 22090 3292
rect 21794 3238 21840 3290
rect 21840 3238 21850 3290
rect 21874 3238 21904 3290
rect 21904 3238 21916 3290
rect 21916 3238 21930 3290
rect 21954 3238 21968 3290
rect 21968 3238 21980 3290
rect 21980 3238 22010 3290
rect 22034 3238 22044 3290
rect 22044 3238 22090 3290
rect 21794 3236 21850 3238
rect 21874 3236 21930 3238
rect 21954 3236 22010 3238
rect 22034 3236 22090 3238
rect 28740 3290 28796 3292
rect 28820 3290 28876 3292
rect 28900 3290 28956 3292
rect 28980 3290 29036 3292
rect 28740 3238 28786 3290
rect 28786 3238 28796 3290
rect 28820 3238 28850 3290
rect 28850 3238 28862 3290
rect 28862 3238 28876 3290
rect 28900 3238 28914 3290
rect 28914 3238 28926 3290
rect 28926 3238 28956 3290
rect 28980 3238 28990 3290
rect 28990 3238 29036 3290
rect 28740 3236 28796 3238
rect 28820 3236 28876 3238
rect 28900 3236 28956 3238
rect 28980 3236 29036 3238
rect 1582 3032 1638 3088
rect 4429 2746 4485 2748
rect 4509 2746 4565 2748
rect 4589 2746 4645 2748
rect 4669 2746 4725 2748
rect 4429 2694 4475 2746
rect 4475 2694 4485 2746
rect 4509 2694 4539 2746
rect 4539 2694 4551 2746
rect 4551 2694 4565 2746
rect 4589 2694 4603 2746
rect 4603 2694 4615 2746
rect 4615 2694 4645 2746
rect 4669 2694 4679 2746
rect 4679 2694 4725 2746
rect 4429 2692 4485 2694
rect 4509 2692 4565 2694
rect 4589 2692 4645 2694
rect 4669 2692 4725 2694
rect 11375 2746 11431 2748
rect 11455 2746 11511 2748
rect 11535 2746 11591 2748
rect 11615 2746 11671 2748
rect 11375 2694 11421 2746
rect 11421 2694 11431 2746
rect 11455 2694 11485 2746
rect 11485 2694 11497 2746
rect 11497 2694 11511 2746
rect 11535 2694 11549 2746
rect 11549 2694 11561 2746
rect 11561 2694 11591 2746
rect 11615 2694 11625 2746
rect 11625 2694 11671 2746
rect 11375 2692 11431 2694
rect 11455 2692 11511 2694
rect 11535 2692 11591 2694
rect 11615 2692 11671 2694
rect 18321 2746 18377 2748
rect 18401 2746 18457 2748
rect 18481 2746 18537 2748
rect 18561 2746 18617 2748
rect 18321 2694 18367 2746
rect 18367 2694 18377 2746
rect 18401 2694 18431 2746
rect 18431 2694 18443 2746
rect 18443 2694 18457 2746
rect 18481 2694 18495 2746
rect 18495 2694 18507 2746
rect 18507 2694 18537 2746
rect 18561 2694 18571 2746
rect 18571 2694 18617 2746
rect 18321 2692 18377 2694
rect 18401 2692 18457 2694
rect 18481 2692 18537 2694
rect 18561 2692 18617 2694
rect 25267 2746 25323 2748
rect 25347 2746 25403 2748
rect 25427 2746 25483 2748
rect 25507 2746 25563 2748
rect 25267 2694 25313 2746
rect 25313 2694 25323 2746
rect 25347 2694 25377 2746
rect 25377 2694 25389 2746
rect 25389 2694 25403 2746
rect 25427 2694 25441 2746
rect 25441 2694 25453 2746
rect 25453 2694 25483 2746
rect 25507 2694 25517 2746
rect 25517 2694 25563 2746
rect 25267 2692 25323 2694
rect 25347 2692 25403 2694
rect 25427 2692 25483 2694
rect 25507 2692 25563 2694
rect 28354 2624 28410 2680
rect 7902 2202 7958 2204
rect 7982 2202 8038 2204
rect 8062 2202 8118 2204
rect 8142 2202 8198 2204
rect 7902 2150 7948 2202
rect 7948 2150 7958 2202
rect 7982 2150 8012 2202
rect 8012 2150 8024 2202
rect 8024 2150 8038 2202
rect 8062 2150 8076 2202
rect 8076 2150 8088 2202
rect 8088 2150 8118 2202
rect 8142 2150 8152 2202
rect 8152 2150 8198 2202
rect 7902 2148 7958 2150
rect 7982 2148 8038 2150
rect 8062 2148 8118 2150
rect 8142 2148 8198 2150
rect 14848 2202 14904 2204
rect 14928 2202 14984 2204
rect 15008 2202 15064 2204
rect 15088 2202 15144 2204
rect 14848 2150 14894 2202
rect 14894 2150 14904 2202
rect 14928 2150 14958 2202
rect 14958 2150 14970 2202
rect 14970 2150 14984 2202
rect 15008 2150 15022 2202
rect 15022 2150 15034 2202
rect 15034 2150 15064 2202
rect 15088 2150 15098 2202
rect 15098 2150 15144 2202
rect 14848 2148 14904 2150
rect 14928 2148 14984 2150
rect 15008 2148 15064 2150
rect 15088 2148 15144 2150
rect 21794 2202 21850 2204
rect 21874 2202 21930 2204
rect 21954 2202 22010 2204
rect 22034 2202 22090 2204
rect 21794 2150 21840 2202
rect 21840 2150 21850 2202
rect 21874 2150 21904 2202
rect 21904 2150 21916 2202
rect 21916 2150 21930 2202
rect 21954 2150 21968 2202
rect 21968 2150 21980 2202
rect 21980 2150 22010 2202
rect 22034 2150 22044 2202
rect 22044 2150 22090 2202
rect 21794 2148 21850 2150
rect 21874 2148 21930 2150
rect 21954 2148 22010 2150
rect 22034 2148 22090 2150
rect 28740 2202 28796 2204
rect 28820 2202 28876 2204
rect 28900 2202 28956 2204
rect 28980 2202 29036 2204
rect 28740 2150 28786 2202
rect 28786 2150 28796 2202
rect 28820 2150 28850 2202
rect 28850 2150 28862 2202
rect 28862 2150 28876 2202
rect 28900 2150 28914 2202
rect 28914 2150 28926 2202
rect 28926 2150 28956 2202
rect 28980 2150 28990 2202
rect 28990 2150 29036 2202
rect 28740 2148 28796 2150
rect 28820 2148 28876 2150
rect 28900 2148 28956 2150
rect 28980 2148 29036 2150
<< metal3 >>
rect 27705 31922 27771 31925
rect 29200 31922 30000 31952
rect 27705 31920 30000 31922
rect 27705 31864 27710 31920
rect 27766 31864 30000 31920
rect 27705 31862 30000 31864
rect 27705 31859 27771 31862
rect 29200 31832 30000 31862
rect 14549 31786 14615 31789
rect 16430 31786 16436 31788
rect 14549 31784 16436 31786
rect 14549 31728 14554 31784
rect 14610 31728 16436 31784
rect 14549 31726 16436 31728
rect 14549 31723 14615 31726
rect 16430 31724 16436 31726
rect 16500 31724 16506 31788
rect 7892 31584 8208 31585
rect 7892 31520 7898 31584
rect 7962 31520 7978 31584
rect 8042 31520 8058 31584
rect 8122 31520 8138 31584
rect 8202 31520 8208 31584
rect 7892 31519 8208 31520
rect 14838 31584 15154 31585
rect 14838 31520 14844 31584
rect 14908 31520 14924 31584
rect 14988 31520 15004 31584
rect 15068 31520 15084 31584
rect 15148 31520 15154 31584
rect 14838 31519 15154 31520
rect 21784 31584 22100 31585
rect 21784 31520 21790 31584
rect 21854 31520 21870 31584
rect 21934 31520 21950 31584
rect 22014 31520 22030 31584
rect 22094 31520 22100 31584
rect 21784 31519 22100 31520
rect 28730 31584 29046 31585
rect 28730 31520 28736 31584
rect 28800 31520 28816 31584
rect 28880 31520 28896 31584
rect 28960 31520 28976 31584
rect 29040 31520 29046 31584
rect 28730 31519 29046 31520
rect 5441 31378 5507 31381
rect 15326 31378 15332 31380
rect 5441 31376 15332 31378
rect 5441 31320 5446 31376
rect 5502 31320 15332 31376
rect 5441 31318 15332 31320
rect 5441 31315 5507 31318
rect 15326 31316 15332 31318
rect 15396 31316 15402 31380
rect 6637 31242 6703 31245
rect 18689 31242 18755 31245
rect 6637 31240 18755 31242
rect 6637 31184 6642 31240
rect 6698 31184 18694 31240
rect 18750 31184 18755 31240
rect 6637 31182 18755 31184
rect 6637 31179 6703 31182
rect 18689 31179 18755 31182
rect 28349 31242 28415 31245
rect 29200 31242 30000 31272
rect 28349 31240 30000 31242
rect 28349 31184 28354 31240
rect 28410 31184 30000 31240
rect 28349 31182 30000 31184
rect 28349 31179 28415 31182
rect 29200 31152 30000 31182
rect 11789 31106 11855 31109
rect 16665 31106 16731 31109
rect 17861 31106 17927 31109
rect 11789 31104 17927 31106
rect 11789 31048 11794 31104
rect 11850 31048 16670 31104
rect 16726 31048 17866 31104
rect 17922 31048 17927 31104
rect 11789 31046 17927 31048
rect 11789 31043 11855 31046
rect 16665 31043 16731 31046
rect 17861 31043 17927 31046
rect 4419 31040 4735 31041
rect 0 30880 800 31000
rect 4419 30976 4425 31040
rect 4489 30976 4505 31040
rect 4569 30976 4585 31040
rect 4649 30976 4665 31040
rect 4729 30976 4735 31040
rect 4419 30975 4735 30976
rect 11365 31040 11681 31041
rect 11365 30976 11371 31040
rect 11435 30976 11451 31040
rect 11515 30976 11531 31040
rect 11595 30976 11611 31040
rect 11675 30976 11681 31040
rect 11365 30975 11681 30976
rect 18311 31040 18627 31041
rect 18311 30976 18317 31040
rect 18381 30976 18397 31040
rect 18461 30976 18477 31040
rect 18541 30976 18557 31040
rect 18621 30976 18627 31040
rect 18311 30975 18627 30976
rect 25257 31040 25573 31041
rect 25257 30976 25263 31040
rect 25327 30976 25343 31040
rect 25407 30976 25423 31040
rect 25487 30976 25503 31040
rect 25567 30976 25573 31040
rect 25257 30975 25573 30976
rect 12709 30970 12775 30973
rect 15377 30970 15443 30973
rect 12709 30968 15443 30970
rect 12709 30912 12714 30968
rect 12770 30912 15382 30968
rect 15438 30912 15443 30968
rect 12709 30910 15443 30912
rect 12709 30907 12775 30910
rect 15377 30907 15443 30910
rect 7557 30834 7623 30837
rect 19793 30834 19859 30837
rect 7557 30832 19859 30834
rect 7557 30776 7562 30832
rect 7618 30776 19798 30832
rect 19854 30776 19859 30832
rect 7557 30774 19859 30776
rect 7557 30771 7623 30774
rect 19793 30771 19859 30774
rect 7189 30698 7255 30701
rect 11789 30698 11855 30701
rect 7189 30696 11855 30698
rect 7189 30640 7194 30696
rect 7250 30640 11794 30696
rect 11850 30640 11855 30696
rect 7189 30638 11855 30640
rect 7189 30635 7255 30638
rect 11789 30635 11855 30638
rect 12157 30698 12223 30701
rect 14273 30698 14339 30701
rect 16481 30698 16547 30701
rect 12157 30696 14339 30698
rect 12157 30640 12162 30696
rect 12218 30640 14278 30696
rect 14334 30640 14339 30696
rect 12157 30638 14339 30640
rect 12157 30635 12223 30638
rect 14273 30635 14339 30638
rect 14414 30696 16547 30698
rect 14414 30640 16486 30696
rect 16542 30640 16547 30696
rect 14414 30638 16547 30640
rect 11145 30562 11211 30565
rect 14414 30562 14474 30638
rect 16481 30635 16547 30638
rect 11145 30560 14474 30562
rect 11145 30504 11150 30560
rect 11206 30504 14474 30560
rect 11145 30502 14474 30504
rect 11145 30499 11211 30502
rect 7892 30496 8208 30497
rect 7892 30432 7898 30496
rect 7962 30432 7978 30496
rect 8042 30432 8058 30496
rect 8122 30432 8138 30496
rect 8202 30432 8208 30496
rect 7892 30431 8208 30432
rect 14838 30496 15154 30497
rect 14838 30432 14844 30496
rect 14908 30432 14924 30496
rect 14988 30432 15004 30496
rect 15068 30432 15084 30496
rect 15148 30432 15154 30496
rect 14838 30431 15154 30432
rect 21784 30496 22100 30497
rect 21784 30432 21790 30496
rect 21854 30432 21870 30496
rect 21934 30432 21950 30496
rect 22014 30432 22030 30496
rect 22094 30432 22100 30496
rect 21784 30431 22100 30432
rect 28730 30496 29046 30497
rect 28730 30432 28736 30496
rect 28800 30432 28816 30496
rect 28880 30432 28896 30496
rect 28960 30432 28976 30496
rect 29040 30432 29046 30496
rect 29200 30472 30000 30592
rect 28730 30431 29046 30432
rect 6729 30426 6795 30429
rect 6862 30426 6868 30428
rect 6729 30424 6868 30426
rect 6729 30368 6734 30424
rect 6790 30368 6868 30424
rect 6729 30366 6868 30368
rect 6729 30363 6795 30366
rect 6862 30364 6868 30366
rect 6932 30364 6938 30428
rect 13629 30426 13695 30429
rect 14549 30426 14615 30429
rect 13629 30424 14615 30426
rect 13629 30368 13634 30424
rect 13690 30368 14554 30424
rect 14610 30368 14615 30424
rect 13629 30366 14615 30368
rect 13629 30363 13695 30366
rect 14549 30363 14615 30366
rect 15561 30426 15627 30429
rect 16614 30426 16620 30428
rect 15561 30424 16620 30426
rect 15561 30368 15566 30424
rect 15622 30368 16620 30424
rect 15561 30366 16620 30368
rect 15561 30363 15627 30366
rect 16614 30364 16620 30366
rect 16684 30364 16690 30428
rect 19885 30426 19951 30429
rect 16806 30424 19951 30426
rect 16806 30368 19890 30424
rect 19946 30368 19951 30424
rect 16806 30366 19951 30368
rect 0 30290 800 30320
rect 2865 30290 2931 30293
rect 0 30288 2931 30290
rect 0 30232 2870 30288
rect 2926 30232 2931 30288
rect 0 30230 2931 30232
rect 0 30200 800 30230
rect 2865 30227 2931 30230
rect 6085 30290 6151 30293
rect 7005 30290 7071 30293
rect 6085 30288 7071 30290
rect 6085 30232 6090 30288
rect 6146 30232 7010 30288
rect 7066 30232 7071 30288
rect 6085 30230 7071 30232
rect 6085 30227 6151 30230
rect 7005 30227 7071 30230
rect 9673 30290 9739 30293
rect 11789 30290 11855 30293
rect 16573 30290 16639 30293
rect 9673 30288 11855 30290
rect 9673 30232 9678 30288
rect 9734 30232 11794 30288
rect 11850 30232 11855 30288
rect 9673 30230 11855 30232
rect 9673 30227 9739 30230
rect 11789 30227 11855 30230
rect 12390 30288 16639 30290
rect 12390 30232 16578 30288
rect 16634 30232 16639 30288
rect 12390 30230 16639 30232
rect 2313 30154 2379 30157
rect 12390 30154 12450 30230
rect 16573 30227 16639 30230
rect 2313 30152 12450 30154
rect 2313 30096 2318 30152
rect 2374 30096 12450 30152
rect 2313 30094 12450 30096
rect 2313 30091 2379 30094
rect 14590 30092 14596 30156
rect 14660 30154 14666 30156
rect 16806 30154 16866 30366
rect 19885 30363 19951 30366
rect 19609 30154 19675 30157
rect 14660 30094 16866 30154
rect 16990 30152 19675 30154
rect 16990 30096 19614 30152
rect 19670 30096 19675 30152
rect 16990 30094 19675 30096
rect 14660 30092 14666 30094
rect 12433 30018 12499 30021
rect 13077 30018 13143 30021
rect 16990 30018 17050 30094
rect 19609 30091 19675 30094
rect 12433 30016 17050 30018
rect 12433 29960 12438 30016
rect 12494 29960 13082 30016
rect 13138 29960 17050 30016
rect 12433 29958 17050 29960
rect 12433 29955 12499 29958
rect 13077 29955 13143 29958
rect 4419 29952 4735 29953
rect 4419 29888 4425 29952
rect 4489 29888 4505 29952
rect 4569 29888 4585 29952
rect 4649 29888 4665 29952
rect 4729 29888 4735 29952
rect 4419 29887 4735 29888
rect 11365 29952 11681 29953
rect 11365 29888 11371 29952
rect 11435 29888 11451 29952
rect 11515 29888 11531 29952
rect 11595 29888 11611 29952
rect 11675 29888 11681 29952
rect 11365 29887 11681 29888
rect 18311 29952 18627 29953
rect 18311 29888 18317 29952
rect 18381 29888 18397 29952
rect 18461 29888 18477 29952
rect 18541 29888 18557 29952
rect 18621 29888 18627 29952
rect 18311 29887 18627 29888
rect 25257 29952 25573 29953
rect 25257 29888 25263 29952
rect 25327 29888 25343 29952
rect 25407 29888 25423 29952
rect 25487 29888 25503 29952
rect 25567 29888 25573 29952
rect 25257 29887 25573 29888
rect 13169 29882 13235 29885
rect 14641 29882 14707 29885
rect 13169 29880 14707 29882
rect 13169 29824 13174 29880
rect 13230 29824 14646 29880
rect 14702 29824 14707 29880
rect 13169 29822 14707 29824
rect 13169 29819 13235 29822
rect 14641 29819 14707 29822
rect 14825 29882 14891 29885
rect 17125 29882 17191 29885
rect 14825 29880 17191 29882
rect 14825 29824 14830 29880
rect 14886 29824 17130 29880
rect 17186 29824 17191 29880
rect 14825 29822 17191 29824
rect 14825 29819 14891 29822
rect 17125 29819 17191 29822
rect 28349 29882 28415 29885
rect 29200 29882 30000 29912
rect 28349 29880 30000 29882
rect 28349 29824 28354 29880
rect 28410 29824 30000 29880
rect 28349 29822 30000 29824
rect 28349 29819 28415 29822
rect 29200 29792 30000 29822
rect 12065 29746 12131 29749
rect 15009 29746 15075 29749
rect 12065 29744 15075 29746
rect 12065 29688 12070 29744
rect 12126 29688 15014 29744
rect 15070 29688 15075 29744
rect 12065 29686 15075 29688
rect 12065 29683 12131 29686
rect 15009 29683 15075 29686
rect 15326 29684 15332 29748
rect 15396 29746 15402 29748
rect 15469 29746 15535 29749
rect 15396 29744 15535 29746
rect 15396 29688 15474 29744
rect 15530 29688 15535 29744
rect 15396 29686 15535 29688
rect 15396 29684 15402 29686
rect 15469 29683 15535 29686
rect 15694 29684 15700 29748
rect 15764 29746 15770 29748
rect 16205 29746 16271 29749
rect 15764 29744 16271 29746
rect 15764 29688 16210 29744
rect 16266 29688 16271 29744
rect 15764 29686 16271 29688
rect 15764 29684 15770 29686
rect 16205 29683 16271 29686
rect 0 29610 800 29640
rect 2589 29610 2655 29613
rect 12934 29610 12940 29612
rect 0 29550 1594 29610
rect 0 29520 800 29550
rect 1534 29474 1594 29550
rect 2589 29608 12940 29610
rect 2589 29552 2594 29608
rect 2650 29552 12940 29608
rect 2589 29550 12940 29552
rect 2589 29547 2655 29550
rect 12934 29548 12940 29550
rect 13004 29548 13010 29612
rect 15837 29610 15903 29613
rect 14598 29608 15903 29610
rect 14598 29552 15842 29608
rect 15898 29552 15903 29608
rect 14598 29550 15903 29552
rect 14598 29477 14658 29550
rect 2957 29474 3023 29477
rect 1534 29472 3023 29474
rect 1534 29416 2962 29472
rect 3018 29416 3023 29472
rect 1534 29414 3023 29416
rect 14598 29472 14707 29477
rect 14598 29416 14646 29472
rect 14702 29416 14707 29472
rect 14598 29414 14707 29416
rect 15702 29474 15762 29550
rect 15837 29547 15903 29550
rect 17309 29610 17375 29613
rect 18965 29610 19031 29613
rect 17309 29608 19031 29610
rect 17309 29552 17314 29608
rect 17370 29552 18970 29608
rect 19026 29552 19031 29608
rect 17309 29550 19031 29552
rect 17309 29547 17375 29550
rect 18965 29547 19031 29550
rect 16205 29474 16271 29477
rect 16665 29476 16731 29477
rect 15702 29472 16271 29474
rect 15702 29416 16210 29472
rect 16266 29416 16271 29472
rect 15702 29414 16271 29416
rect 2957 29411 3023 29414
rect 14641 29411 14707 29414
rect 16205 29411 16271 29414
rect 16614 29412 16620 29476
rect 16684 29474 16731 29476
rect 16684 29472 16776 29474
rect 16726 29416 16776 29472
rect 16684 29414 16776 29416
rect 16684 29412 16731 29414
rect 16665 29411 16731 29412
rect 7892 29408 8208 29409
rect 7892 29344 7898 29408
rect 7962 29344 7978 29408
rect 8042 29344 8058 29408
rect 8122 29344 8138 29408
rect 8202 29344 8208 29408
rect 7892 29343 8208 29344
rect 14838 29408 15154 29409
rect 14838 29344 14844 29408
rect 14908 29344 14924 29408
rect 14988 29344 15004 29408
rect 15068 29344 15084 29408
rect 15148 29344 15154 29408
rect 14838 29343 15154 29344
rect 21784 29408 22100 29409
rect 21784 29344 21790 29408
rect 21854 29344 21870 29408
rect 21934 29344 21950 29408
rect 22014 29344 22030 29408
rect 22094 29344 22100 29408
rect 21784 29343 22100 29344
rect 28730 29408 29046 29409
rect 28730 29344 28736 29408
rect 28800 29344 28816 29408
rect 28880 29344 28896 29408
rect 28960 29344 28976 29408
rect 29040 29344 29046 29408
rect 28730 29343 29046 29344
rect 10225 29338 10291 29341
rect 15377 29338 15443 29341
rect 19057 29338 19123 29341
rect 10225 29336 14474 29338
rect 10225 29280 10230 29336
rect 10286 29280 14474 29336
rect 10225 29278 14474 29280
rect 10225 29275 10291 29278
rect 5993 29202 6059 29205
rect 11145 29202 11211 29205
rect 14181 29202 14247 29205
rect 5993 29200 14247 29202
rect 5993 29144 5998 29200
rect 6054 29144 11150 29200
rect 11206 29144 14186 29200
rect 14242 29144 14247 29200
rect 5993 29142 14247 29144
rect 14414 29202 14474 29278
rect 15377 29336 19123 29338
rect 15377 29280 15382 29336
rect 15438 29280 19062 29336
rect 19118 29280 19123 29336
rect 15377 29278 19123 29280
rect 15377 29275 15443 29278
rect 19057 29275 19123 29278
rect 15694 29202 15700 29204
rect 14414 29142 15700 29202
rect 5993 29139 6059 29142
rect 11145 29139 11211 29142
rect 14181 29139 14247 29142
rect 15694 29140 15700 29142
rect 15764 29140 15770 29204
rect 16430 29140 16436 29204
rect 16500 29202 16506 29204
rect 16665 29202 16731 29205
rect 16500 29200 16731 29202
rect 16500 29144 16670 29200
rect 16726 29144 16731 29200
rect 16500 29142 16731 29144
rect 16500 29140 16506 29142
rect 16665 29139 16731 29142
rect 28349 29202 28415 29205
rect 29200 29202 30000 29232
rect 28349 29200 30000 29202
rect 28349 29144 28354 29200
rect 28410 29144 30000 29200
rect 28349 29142 30000 29144
rect 28349 29139 28415 29142
rect 29200 29112 30000 29142
rect 7557 29066 7623 29069
rect 8385 29066 8451 29069
rect 7557 29064 8451 29066
rect 7557 29008 7562 29064
rect 7618 29008 8390 29064
rect 8446 29008 8451 29064
rect 7557 29006 8451 29008
rect 7557 29003 7623 29006
rect 8385 29003 8451 29006
rect 8937 29066 9003 29069
rect 14733 29066 14799 29069
rect 17033 29066 17099 29069
rect 8937 29064 17099 29066
rect 8937 29008 8942 29064
rect 8998 29008 14738 29064
rect 14794 29008 17038 29064
rect 17094 29008 17099 29064
rect 8937 29006 17099 29008
rect 8937 29003 9003 29006
rect 14733 29003 14799 29006
rect 17033 29003 17099 29006
rect 0 28840 800 28960
rect 7097 28930 7163 28933
rect 9857 28930 9923 28933
rect 7097 28928 9923 28930
rect 7097 28872 7102 28928
rect 7158 28872 9862 28928
rect 9918 28872 9923 28928
rect 7097 28870 9923 28872
rect 7097 28867 7163 28870
rect 9857 28867 9923 28870
rect 12249 28930 12315 28933
rect 12709 28930 12775 28933
rect 12249 28928 12775 28930
rect 12249 28872 12254 28928
rect 12310 28872 12714 28928
rect 12770 28872 12775 28928
rect 12249 28870 12775 28872
rect 12249 28867 12315 28870
rect 12709 28867 12775 28870
rect 12893 28930 12959 28933
rect 16757 28930 16823 28933
rect 12893 28928 16823 28930
rect 12893 28872 12898 28928
rect 12954 28872 16762 28928
rect 16818 28872 16823 28928
rect 12893 28870 16823 28872
rect 12893 28867 12959 28870
rect 16757 28867 16823 28870
rect 4419 28864 4735 28865
rect 4419 28800 4425 28864
rect 4489 28800 4505 28864
rect 4569 28800 4585 28864
rect 4649 28800 4665 28864
rect 4729 28800 4735 28864
rect 4419 28799 4735 28800
rect 11365 28864 11681 28865
rect 11365 28800 11371 28864
rect 11435 28800 11451 28864
rect 11515 28800 11531 28864
rect 11595 28800 11611 28864
rect 11675 28800 11681 28864
rect 11365 28799 11681 28800
rect 18311 28864 18627 28865
rect 18311 28800 18317 28864
rect 18381 28800 18397 28864
rect 18461 28800 18477 28864
rect 18541 28800 18557 28864
rect 18621 28800 18627 28864
rect 18311 28799 18627 28800
rect 25257 28864 25573 28865
rect 25257 28800 25263 28864
rect 25327 28800 25343 28864
rect 25407 28800 25423 28864
rect 25487 28800 25503 28864
rect 25567 28800 25573 28864
rect 25257 28799 25573 28800
rect 11789 28794 11855 28797
rect 18137 28794 18203 28797
rect 11789 28792 18203 28794
rect 11789 28736 11794 28792
rect 11850 28736 18142 28792
rect 18198 28736 18203 28792
rect 11789 28734 18203 28736
rect 11789 28731 11855 28734
rect 18137 28731 18203 28734
rect 3233 28658 3299 28661
rect 3969 28658 4035 28661
rect 4153 28658 4219 28661
rect 8661 28658 8727 28661
rect 3233 28656 8727 28658
rect 3233 28600 3238 28656
rect 3294 28600 3974 28656
rect 4030 28600 4158 28656
rect 4214 28600 8666 28656
rect 8722 28600 8727 28656
rect 3233 28598 8727 28600
rect 3233 28595 3299 28598
rect 3969 28595 4035 28598
rect 4153 28595 4219 28598
rect 8661 28595 8727 28598
rect 11789 28658 11855 28661
rect 14089 28658 14155 28661
rect 11789 28656 14155 28658
rect 11789 28600 11794 28656
rect 11850 28600 14094 28656
rect 14150 28600 14155 28656
rect 11789 28598 14155 28600
rect 11789 28595 11855 28598
rect 14089 28595 14155 28598
rect 13169 28522 13235 28525
rect 13905 28522 13971 28525
rect 13169 28520 13971 28522
rect 13169 28464 13174 28520
rect 13230 28464 13910 28520
rect 13966 28464 13971 28520
rect 13169 28462 13971 28464
rect 13169 28459 13235 28462
rect 13905 28459 13971 28462
rect 29200 28432 30000 28552
rect 7892 28320 8208 28321
rect 0 28250 800 28280
rect 7892 28256 7898 28320
rect 7962 28256 7978 28320
rect 8042 28256 8058 28320
rect 8122 28256 8138 28320
rect 8202 28256 8208 28320
rect 7892 28255 8208 28256
rect 14838 28320 15154 28321
rect 14838 28256 14844 28320
rect 14908 28256 14924 28320
rect 14988 28256 15004 28320
rect 15068 28256 15084 28320
rect 15148 28256 15154 28320
rect 14838 28255 15154 28256
rect 21784 28320 22100 28321
rect 21784 28256 21790 28320
rect 21854 28256 21870 28320
rect 21934 28256 21950 28320
rect 22014 28256 22030 28320
rect 22094 28256 22100 28320
rect 21784 28255 22100 28256
rect 28730 28320 29046 28321
rect 28730 28256 28736 28320
rect 28800 28256 28816 28320
rect 28880 28256 28896 28320
rect 28960 28256 28976 28320
rect 29040 28256 29046 28320
rect 28730 28255 29046 28256
rect 1669 28250 1735 28253
rect 0 28248 1735 28250
rect 0 28192 1674 28248
rect 1730 28192 1735 28248
rect 0 28190 1735 28192
rect 0 28160 800 28190
rect 1669 28187 1735 28190
rect 9949 28250 10015 28253
rect 13353 28250 13419 28253
rect 9949 28248 13419 28250
rect 9949 28192 9954 28248
rect 10010 28192 13358 28248
rect 13414 28192 13419 28248
rect 9949 28190 13419 28192
rect 9949 28187 10015 28190
rect 13353 28187 13419 28190
rect 9673 28114 9739 28117
rect 15009 28114 15075 28117
rect 9673 28112 15075 28114
rect 9673 28056 9678 28112
rect 9734 28056 15014 28112
rect 15070 28056 15075 28112
rect 9673 28054 15075 28056
rect 9673 28051 9739 28054
rect 15009 28051 15075 28054
rect 2037 27978 2103 27981
rect 12617 27978 12683 27981
rect 12750 27978 12756 27980
rect 2037 27976 12450 27978
rect 2037 27920 2042 27976
rect 2098 27920 12450 27976
rect 2037 27918 12450 27920
rect 2037 27915 2103 27918
rect 4419 27776 4735 27777
rect 4419 27712 4425 27776
rect 4489 27712 4505 27776
rect 4569 27712 4585 27776
rect 4649 27712 4665 27776
rect 4729 27712 4735 27776
rect 4419 27711 4735 27712
rect 11365 27776 11681 27777
rect 11365 27712 11371 27776
rect 11435 27712 11451 27776
rect 11515 27712 11531 27776
rect 11595 27712 11611 27776
rect 11675 27712 11681 27776
rect 11365 27711 11681 27712
rect 12390 27706 12450 27918
rect 12617 27976 12756 27978
rect 12617 27920 12622 27976
rect 12678 27920 12756 27976
rect 12617 27918 12756 27920
rect 12617 27915 12683 27918
rect 12750 27916 12756 27918
rect 12820 27916 12826 27980
rect 13445 27978 13511 27981
rect 15469 27978 15535 27981
rect 13445 27976 15535 27978
rect 13445 27920 13450 27976
rect 13506 27920 15474 27976
rect 15530 27920 15535 27976
rect 13445 27918 15535 27920
rect 13445 27915 13511 27918
rect 15469 27915 15535 27918
rect 12617 27842 12683 27845
rect 17953 27842 18019 27845
rect 12617 27840 18019 27842
rect 12617 27784 12622 27840
rect 12678 27784 17958 27840
rect 18014 27784 18019 27840
rect 12617 27782 18019 27784
rect 12617 27779 12683 27782
rect 17953 27779 18019 27782
rect 28349 27842 28415 27845
rect 29200 27842 30000 27872
rect 28349 27840 30000 27842
rect 28349 27784 28354 27840
rect 28410 27784 30000 27840
rect 28349 27782 30000 27784
rect 28349 27779 28415 27782
rect 18311 27776 18627 27777
rect 18311 27712 18317 27776
rect 18381 27712 18397 27776
rect 18461 27712 18477 27776
rect 18541 27712 18557 27776
rect 18621 27712 18627 27776
rect 18311 27711 18627 27712
rect 25257 27776 25573 27777
rect 25257 27712 25263 27776
rect 25327 27712 25343 27776
rect 25407 27712 25423 27776
rect 25487 27712 25503 27776
rect 25567 27712 25573 27776
rect 29200 27752 30000 27782
rect 25257 27711 25573 27712
rect 13813 27706 13879 27709
rect 14181 27706 14247 27709
rect 17125 27706 17191 27709
rect 12390 27646 13738 27706
rect 0 27570 800 27600
rect 2773 27570 2839 27573
rect 0 27568 2839 27570
rect 0 27512 2778 27568
rect 2834 27512 2839 27568
rect 0 27510 2839 27512
rect 0 27480 800 27510
rect 2773 27507 2839 27510
rect 10961 27570 11027 27573
rect 13678 27570 13738 27646
rect 13813 27704 17191 27706
rect 13813 27648 13818 27704
rect 13874 27648 14186 27704
rect 14242 27648 17130 27704
rect 17186 27648 17191 27704
rect 13813 27646 17191 27648
rect 13813 27643 13879 27646
rect 14181 27643 14247 27646
rect 17125 27643 17191 27646
rect 15929 27570 15995 27573
rect 10961 27568 13370 27570
rect 10961 27512 10966 27568
rect 11022 27512 13370 27568
rect 10961 27510 13370 27512
rect 13678 27568 15995 27570
rect 13678 27512 15934 27568
rect 15990 27512 15995 27568
rect 13678 27510 15995 27512
rect 10961 27507 11027 27510
rect 2221 27434 2287 27437
rect 6453 27434 6519 27437
rect 2221 27432 6519 27434
rect 2221 27376 2226 27432
rect 2282 27376 6458 27432
rect 6514 27376 6519 27432
rect 2221 27374 6519 27376
rect 2221 27371 2287 27374
rect 6453 27371 6519 27374
rect 6862 27372 6868 27436
rect 6932 27434 6938 27436
rect 8753 27434 8819 27437
rect 13169 27434 13235 27437
rect 6932 27374 8586 27434
rect 6932 27372 6938 27374
rect 7892 27232 8208 27233
rect 7892 27168 7898 27232
rect 7962 27168 7978 27232
rect 8042 27168 8058 27232
rect 8122 27168 8138 27232
rect 8202 27168 8208 27232
rect 7892 27167 8208 27168
rect 4705 27162 4771 27165
rect 6269 27162 6335 27165
rect 4705 27160 6335 27162
rect 4705 27104 4710 27160
rect 4766 27104 6274 27160
rect 6330 27104 6335 27160
rect 4705 27102 6335 27104
rect 8526 27162 8586 27374
rect 8753 27432 13235 27434
rect 8753 27376 8758 27432
rect 8814 27376 13174 27432
rect 13230 27376 13235 27432
rect 8753 27374 13235 27376
rect 13310 27434 13370 27510
rect 15929 27507 15995 27510
rect 13905 27434 13971 27437
rect 15653 27434 15719 27437
rect 13310 27432 13971 27434
rect 13310 27376 13910 27432
rect 13966 27376 13971 27432
rect 13310 27374 13971 27376
rect 8753 27371 8819 27374
rect 13169 27371 13235 27374
rect 13905 27371 13971 27374
rect 14046 27432 15719 27434
rect 14046 27376 15658 27432
rect 15714 27376 15719 27432
rect 14046 27374 15719 27376
rect 12985 27300 13051 27301
rect 12934 27236 12940 27300
rect 13004 27298 13051 27300
rect 13445 27298 13511 27301
rect 14046 27298 14106 27374
rect 15653 27371 15719 27374
rect 28349 27434 28415 27437
rect 28349 27432 29378 27434
rect 28349 27376 28354 27432
rect 28410 27376 29378 27432
rect 28349 27374 29378 27376
rect 28349 27371 28415 27374
rect 13004 27296 13096 27298
rect 13046 27240 13096 27296
rect 13004 27238 13096 27240
rect 13445 27296 14106 27298
rect 13445 27240 13450 27296
rect 13506 27240 14106 27296
rect 13445 27238 14106 27240
rect 13004 27236 13051 27238
rect 12985 27235 13051 27236
rect 13445 27235 13511 27238
rect 14838 27232 15154 27233
rect 14838 27168 14844 27232
rect 14908 27168 14924 27232
rect 14988 27168 15004 27232
rect 15068 27168 15084 27232
rect 15148 27168 15154 27232
rect 14838 27167 15154 27168
rect 21784 27232 22100 27233
rect 21784 27168 21790 27232
rect 21854 27168 21870 27232
rect 21934 27168 21950 27232
rect 22014 27168 22030 27232
rect 22094 27168 22100 27232
rect 21784 27167 22100 27168
rect 28730 27232 29046 27233
rect 28730 27168 28736 27232
rect 28800 27168 28816 27232
rect 28880 27168 28896 27232
rect 28960 27168 28976 27232
rect 29040 27168 29046 27232
rect 29318 27192 29378 27374
rect 28730 27167 29046 27168
rect 12433 27162 12499 27165
rect 12985 27162 13051 27165
rect 8526 27102 9690 27162
rect 4705 27099 4771 27102
rect 6269 27099 6335 27102
rect 3233 27026 3299 27029
rect 9029 27026 9095 27029
rect 3233 27024 9095 27026
rect 3233 26968 3238 27024
rect 3294 26968 9034 27024
rect 9090 26968 9095 27024
rect 3233 26966 9095 26968
rect 9630 27026 9690 27102
rect 12433 27160 13051 27162
rect 12433 27104 12438 27160
rect 12494 27104 12990 27160
rect 13046 27104 13051 27160
rect 12433 27102 13051 27104
rect 12433 27099 12499 27102
rect 12985 27099 13051 27102
rect 29200 27072 30000 27192
rect 13169 27026 13235 27029
rect 9630 27024 13235 27026
rect 9630 26968 13174 27024
rect 13230 26968 13235 27024
rect 9630 26966 13235 26968
rect 3233 26963 3299 26966
rect 9029 26963 9095 26966
rect 13169 26963 13235 26966
rect 14089 27026 14155 27029
rect 15745 27026 15811 27029
rect 14089 27024 15811 27026
rect 14089 26968 14094 27024
rect 14150 26968 15750 27024
rect 15806 26968 15811 27024
rect 14089 26966 15811 26968
rect 14089 26963 14155 26966
rect 15745 26963 15811 26966
rect 0 26800 800 26920
rect 3693 26890 3759 26893
rect 13445 26890 13511 26893
rect 3693 26888 13511 26890
rect 3693 26832 3698 26888
rect 3754 26832 13450 26888
rect 13506 26832 13511 26888
rect 3693 26830 13511 26832
rect 3693 26827 3759 26830
rect 13445 26827 13511 26830
rect 5717 26754 5783 26757
rect 6361 26754 6427 26757
rect 5717 26752 6427 26754
rect 5717 26696 5722 26752
rect 5778 26696 6366 26752
rect 6422 26696 6427 26752
rect 5717 26694 6427 26696
rect 5717 26691 5783 26694
rect 6361 26691 6427 26694
rect 12525 26754 12591 26757
rect 14457 26754 14523 26757
rect 17309 26754 17375 26757
rect 12525 26752 17375 26754
rect 12525 26696 12530 26752
rect 12586 26696 14462 26752
rect 14518 26696 17314 26752
rect 17370 26696 17375 26752
rect 12525 26694 17375 26696
rect 12525 26691 12591 26694
rect 14457 26691 14523 26694
rect 17309 26691 17375 26694
rect 4419 26688 4735 26689
rect 4419 26624 4425 26688
rect 4489 26624 4505 26688
rect 4569 26624 4585 26688
rect 4649 26624 4665 26688
rect 4729 26624 4735 26688
rect 4419 26623 4735 26624
rect 11365 26688 11681 26689
rect 11365 26624 11371 26688
rect 11435 26624 11451 26688
rect 11515 26624 11531 26688
rect 11595 26624 11611 26688
rect 11675 26624 11681 26688
rect 11365 26623 11681 26624
rect 18311 26688 18627 26689
rect 18311 26624 18317 26688
rect 18381 26624 18397 26688
rect 18461 26624 18477 26688
rect 18541 26624 18557 26688
rect 18621 26624 18627 26688
rect 18311 26623 18627 26624
rect 25257 26688 25573 26689
rect 25257 26624 25263 26688
rect 25327 26624 25343 26688
rect 25407 26624 25423 26688
rect 25487 26624 25503 26688
rect 25567 26624 25573 26688
rect 25257 26623 25573 26624
rect 6637 26618 6703 26621
rect 7649 26618 7715 26621
rect 8753 26618 8819 26621
rect 17493 26618 17559 26621
rect 6637 26616 7715 26618
rect 6637 26560 6642 26616
rect 6698 26560 7654 26616
rect 7710 26560 7715 26616
rect 6637 26558 7715 26560
rect 6637 26555 6703 26558
rect 7649 26555 7715 26558
rect 7790 26616 8819 26618
rect 7790 26560 8758 26616
rect 8814 26560 8819 26616
rect 7790 26558 8819 26560
rect 4429 26482 4495 26485
rect 7790 26482 7850 26558
rect 8753 26555 8819 26558
rect 12390 26616 17559 26618
rect 12390 26560 17498 26616
rect 17554 26560 17559 26616
rect 12390 26558 17559 26560
rect 4429 26480 7850 26482
rect 4429 26424 4434 26480
rect 4490 26424 7850 26480
rect 4429 26422 7850 26424
rect 8385 26482 8451 26485
rect 12390 26482 12450 26558
rect 17493 26555 17559 26558
rect 8385 26480 12450 26482
rect 8385 26424 8390 26480
rect 8446 26424 12450 26480
rect 8385 26422 12450 26424
rect 13629 26482 13695 26485
rect 14590 26482 14596 26484
rect 13629 26480 14596 26482
rect 13629 26424 13634 26480
rect 13690 26424 14596 26480
rect 13629 26422 14596 26424
rect 4429 26419 4495 26422
rect 8385 26419 8451 26422
rect 13629 26419 13695 26422
rect 14590 26420 14596 26422
rect 14660 26420 14666 26484
rect 29200 26392 30000 26512
rect 2589 26346 2655 26349
rect 5533 26346 5599 26349
rect 2589 26344 5599 26346
rect 2589 26288 2594 26344
rect 2650 26288 5538 26344
rect 5594 26288 5599 26344
rect 2589 26286 5599 26288
rect 2589 26283 2655 26286
rect 5533 26283 5599 26286
rect 12433 26346 12499 26349
rect 14089 26346 14155 26349
rect 16297 26346 16363 26349
rect 12433 26344 14155 26346
rect 12433 26288 12438 26344
rect 12494 26288 14094 26344
rect 14150 26288 14155 26344
rect 12433 26286 14155 26288
rect 12433 26283 12499 26286
rect 14089 26283 14155 26286
rect 14230 26344 16363 26346
rect 14230 26288 16302 26344
rect 16358 26288 16363 26344
rect 14230 26286 16363 26288
rect 0 26210 800 26240
rect 1577 26210 1643 26213
rect 0 26208 1643 26210
rect 0 26152 1582 26208
rect 1638 26152 1643 26208
rect 0 26150 1643 26152
rect 0 26120 800 26150
rect 1577 26147 1643 26150
rect 2313 26210 2379 26213
rect 5993 26210 6059 26213
rect 2313 26208 6059 26210
rect 2313 26152 2318 26208
rect 2374 26152 5998 26208
rect 6054 26152 6059 26208
rect 2313 26150 6059 26152
rect 2313 26147 2379 26150
rect 5993 26147 6059 26150
rect 10317 26210 10383 26213
rect 14230 26210 14290 26286
rect 16297 26283 16363 26286
rect 10317 26208 14290 26210
rect 10317 26152 10322 26208
rect 10378 26152 14290 26208
rect 10317 26150 14290 26152
rect 10317 26147 10383 26150
rect 7892 26144 8208 26145
rect 7892 26080 7898 26144
rect 7962 26080 7978 26144
rect 8042 26080 8058 26144
rect 8122 26080 8138 26144
rect 8202 26080 8208 26144
rect 7892 26079 8208 26080
rect 14838 26144 15154 26145
rect 14838 26080 14844 26144
rect 14908 26080 14924 26144
rect 14988 26080 15004 26144
rect 15068 26080 15084 26144
rect 15148 26080 15154 26144
rect 14838 26079 15154 26080
rect 21784 26144 22100 26145
rect 21784 26080 21790 26144
rect 21854 26080 21870 26144
rect 21934 26080 21950 26144
rect 22014 26080 22030 26144
rect 22094 26080 22100 26144
rect 21784 26079 22100 26080
rect 28730 26144 29046 26145
rect 28730 26080 28736 26144
rect 28800 26080 28816 26144
rect 28880 26080 28896 26144
rect 28960 26080 28976 26144
rect 29040 26080 29046 26144
rect 28730 26079 29046 26080
rect 3785 26074 3851 26077
rect 7189 26074 7255 26077
rect 3785 26072 7255 26074
rect 3785 26016 3790 26072
rect 3846 26016 7194 26072
rect 7250 26016 7255 26072
rect 3785 26014 7255 26016
rect 3785 26011 3851 26014
rect 7189 26011 7255 26014
rect 9857 26074 9923 26077
rect 10409 26074 10475 26077
rect 12985 26074 13051 26077
rect 9857 26072 13051 26074
rect 9857 26016 9862 26072
rect 9918 26016 10414 26072
rect 10470 26016 12990 26072
rect 13046 26016 13051 26072
rect 9857 26014 13051 26016
rect 9857 26011 9923 26014
rect 10409 26011 10475 26014
rect 12985 26011 13051 26014
rect 5257 25938 5323 25941
rect 11697 25938 11763 25941
rect 5257 25936 11763 25938
rect 5257 25880 5262 25936
rect 5318 25880 11702 25936
rect 11758 25880 11763 25936
rect 5257 25878 11763 25880
rect 5257 25875 5323 25878
rect 11697 25875 11763 25878
rect 11973 25938 12039 25941
rect 16021 25938 16087 25941
rect 11973 25936 16087 25938
rect 11973 25880 11978 25936
rect 12034 25880 16026 25936
rect 16082 25880 16087 25936
rect 11973 25878 16087 25880
rect 11973 25875 12039 25878
rect 16021 25875 16087 25878
rect 3233 25802 3299 25805
rect 12617 25802 12683 25805
rect 3233 25800 12683 25802
rect 3233 25744 3238 25800
rect 3294 25744 12622 25800
rect 12678 25744 12683 25800
rect 3233 25742 12683 25744
rect 3233 25739 3299 25742
rect 12617 25739 12683 25742
rect 28349 25802 28415 25805
rect 29200 25802 30000 25832
rect 28349 25800 30000 25802
rect 28349 25744 28354 25800
rect 28410 25744 30000 25800
rect 28349 25742 30000 25744
rect 28349 25739 28415 25742
rect 29200 25712 30000 25742
rect 4419 25600 4735 25601
rect 0 25530 800 25560
rect 4419 25536 4425 25600
rect 4489 25536 4505 25600
rect 4569 25536 4585 25600
rect 4649 25536 4665 25600
rect 4729 25536 4735 25600
rect 4419 25535 4735 25536
rect 11365 25600 11681 25601
rect 11365 25536 11371 25600
rect 11435 25536 11451 25600
rect 11515 25536 11531 25600
rect 11595 25536 11611 25600
rect 11675 25536 11681 25600
rect 11365 25535 11681 25536
rect 18311 25600 18627 25601
rect 18311 25536 18317 25600
rect 18381 25536 18397 25600
rect 18461 25536 18477 25600
rect 18541 25536 18557 25600
rect 18621 25536 18627 25600
rect 18311 25535 18627 25536
rect 25257 25600 25573 25601
rect 25257 25536 25263 25600
rect 25327 25536 25343 25600
rect 25407 25536 25423 25600
rect 25487 25536 25503 25600
rect 25567 25536 25573 25600
rect 25257 25535 25573 25536
rect 2313 25530 2379 25533
rect 0 25528 2379 25530
rect 0 25472 2318 25528
rect 2374 25472 2379 25528
rect 0 25470 2379 25472
rect 0 25440 800 25470
rect 2313 25467 2379 25470
rect 6453 25530 6519 25533
rect 7557 25530 7623 25533
rect 6453 25528 7623 25530
rect 6453 25472 6458 25528
rect 6514 25472 7562 25528
rect 7618 25472 7623 25528
rect 6453 25470 7623 25472
rect 6453 25467 6519 25470
rect 7557 25467 7623 25470
rect 7465 25394 7531 25397
rect 7833 25394 7899 25397
rect 7465 25392 7899 25394
rect 7465 25336 7470 25392
rect 7526 25336 7838 25392
rect 7894 25336 7899 25392
rect 7465 25334 7899 25336
rect 7465 25331 7531 25334
rect 7833 25331 7899 25334
rect 9765 25394 9831 25397
rect 11053 25394 11119 25397
rect 9765 25392 11119 25394
rect 9765 25336 9770 25392
rect 9826 25336 11058 25392
rect 11114 25336 11119 25392
rect 9765 25334 11119 25336
rect 9765 25331 9831 25334
rect 11053 25331 11119 25334
rect 28349 25394 28415 25397
rect 28349 25392 29378 25394
rect 28349 25336 28354 25392
rect 28410 25336 29378 25392
rect 28349 25334 29378 25336
rect 28349 25331 28415 25334
rect 4245 25258 4311 25261
rect 10593 25258 10659 25261
rect 4245 25256 10659 25258
rect 4245 25200 4250 25256
rect 4306 25200 10598 25256
rect 10654 25200 10659 25256
rect 4245 25198 10659 25200
rect 4245 25195 4311 25198
rect 10593 25195 10659 25198
rect 29318 25152 29378 25334
rect 7892 25056 8208 25057
rect 7892 24992 7898 25056
rect 7962 24992 7978 25056
rect 8042 24992 8058 25056
rect 8122 24992 8138 25056
rect 8202 24992 8208 25056
rect 7892 24991 8208 24992
rect 14838 25056 15154 25057
rect 14838 24992 14844 25056
rect 14908 24992 14924 25056
rect 14988 24992 15004 25056
rect 15068 24992 15084 25056
rect 15148 24992 15154 25056
rect 14838 24991 15154 24992
rect 21784 25056 22100 25057
rect 21784 24992 21790 25056
rect 21854 24992 21870 25056
rect 21934 24992 21950 25056
rect 22014 24992 22030 25056
rect 22094 24992 22100 25056
rect 21784 24991 22100 24992
rect 28730 25056 29046 25057
rect 28730 24992 28736 25056
rect 28800 24992 28816 25056
rect 28880 24992 28896 25056
rect 28960 24992 28976 25056
rect 29040 24992 29046 25056
rect 29200 25032 30000 25152
rect 28730 24991 29046 24992
rect 5165 24986 5231 24989
rect 7557 24986 7623 24989
rect 5165 24984 7623 24986
rect 5165 24928 5170 24984
rect 5226 24928 7562 24984
rect 7618 24928 7623 24984
rect 5165 24926 7623 24928
rect 5165 24923 5231 24926
rect 7557 24923 7623 24926
rect 0 24760 800 24880
rect 3325 24850 3391 24853
rect 11697 24850 11763 24853
rect 3325 24848 11763 24850
rect 3325 24792 3330 24848
rect 3386 24792 11702 24848
rect 11758 24792 11763 24848
rect 3325 24790 11763 24792
rect 3325 24787 3391 24790
rect 11697 24787 11763 24790
rect 8661 24714 8727 24717
rect 9581 24714 9647 24717
rect 8661 24712 9647 24714
rect 8661 24656 8666 24712
rect 8722 24656 9586 24712
rect 9642 24656 9647 24712
rect 8661 24654 9647 24656
rect 8661 24651 8727 24654
rect 9581 24651 9647 24654
rect 4419 24512 4735 24513
rect 4419 24448 4425 24512
rect 4489 24448 4505 24512
rect 4569 24448 4585 24512
rect 4649 24448 4665 24512
rect 4729 24448 4735 24512
rect 4419 24447 4735 24448
rect 11365 24512 11681 24513
rect 11365 24448 11371 24512
rect 11435 24448 11451 24512
rect 11515 24448 11531 24512
rect 11595 24448 11611 24512
rect 11675 24448 11681 24512
rect 11365 24447 11681 24448
rect 18311 24512 18627 24513
rect 18311 24448 18317 24512
rect 18381 24448 18397 24512
rect 18461 24448 18477 24512
rect 18541 24448 18557 24512
rect 18621 24448 18627 24512
rect 18311 24447 18627 24448
rect 25257 24512 25573 24513
rect 25257 24448 25263 24512
rect 25327 24448 25343 24512
rect 25407 24448 25423 24512
rect 25487 24448 25503 24512
rect 25567 24448 25573 24512
rect 25257 24447 25573 24448
rect 29200 24352 30000 24472
rect 0 24170 800 24200
rect 1577 24170 1643 24173
rect 0 24168 1643 24170
rect 0 24112 1582 24168
rect 1638 24112 1643 24168
rect 0 24110 1643 24112
rect 0 24080 800 24110
rect 1577 24107 1643 24110
rect 7892 23968 8208 23969
rect 7892 23904 7898 23968
rect 7962 23904 7978 23968
rect 8042 23904 8058 23968
rect 8122 23904 8138 23968
rect 8202 23904 8208 23968
rect 7892 23903 8208 23904
rect 14838 23968 15154 23969
rect 14838 23904 14844 23968
rect 14908 23904 14924 23968
rect 14988 23904 15004 23968
rect 15068 23904 15084 23968
rect 15148 23904 15154 23968
rect 14838 23903 15154 23904
rect 21784 23968 22100 23969
rect 21784 23904 21790 23968
rect 21854 23904 21870 23968
rect 21934 23904 21950 23968
rect 22014 23904 22030 23968
rect 22094 23904 22100 23968
rect 21784 23903 22100 23904
rect 28730 23968 29046 23969
rect 28730 23904 28736 23968
rect 28800 23904 28816 23968
rect 28880 23904 28896 23968
rect 28960 23904 28976 23968
rect 29040 23904 29046 23968
rect 28730 23903 29046 23904
rect 28349 23762 28415 23765
rect 29200 23762 30000 23792
rect 28349 23760 30000 23762
rect 28349 23704 28354 23760
rect 28410 23704 30000 23760
rect 28349 23702 30000 23704
rect 28349 23699 28415 23702
rect 29200 23672 30000 23702
rect 0 23490 800 23520
rect 1577 23490 1643 23493
rect 0 23488 1643 23490
rect 0 23432 1582 23488
rect 1638 23432 1643 23488
rect 0 23430 1643 23432
rect 0 23400 800 23430
rect 1577 23427 1643 23430
rect 4419 23424 4735 23425
rect 4419 23360 4425 23424
rect 4489 23360 4505 23424
rect 4569 23360 4585 23424
rect 4649 23360 4665 23424
rect 4729 23360 4735 23424
rect 4419 23359 4735 23360
rect 11365 23424 11681 23425
rect 11365 23360 11371 23424
rect 11435 23360 11451 23424
rect 11515 23360 11531 23424
rect 11595 23360 11611 23424
rect 11675 23360 11681 23424
rect 11365 23359 11681 23360
rect 18311 23424 18627 23425
rect 18311 23360 18317 23424
rect 18381 23360 18397 23424
rect 18461 23360 18477 23424
rect 18541 23360 18557 23424
rect 18621 23360 18627 23424
rect 18311 23359 18627 23360
rect 25257 23424 25573 23425
rect 25257 23360 25263 23424
rect 25327 23360 25343 23424
rect 25407 23360 25423 23424
rect 25487 23360 25503 23424
rect 25567 23360 25573 23424
rect 25257 23359 25573 23360
rect 28349 23082 28415 23085
rect 29200 23082 30000 23112
rect 28349 23080 30000 23082
rect 28349 23024 28354 23080
rect 28410 23024 30000 23080
rect 28349 23022 30000 23024
rect 28349 23019 28415 23022
rect 29200 22992 30000 23022
rect 7892 22880 8208 22881
rect 0 22720 800 22840
rect 7892 22816 7898 22880
rect 7962 22816 7978 22880
rect 8042 22816 8058 22880
rect 8122 22816 8138 22880
rect 8202 22816 8208 22880
rect 7892 22815 8208 22816
rect 14838 22880 15154 22881
rect 14838 22816 14844 22880
rect 14908 22816 14924 22880
rect 14988 22816 15004 22880
rect 15068 22816 15084 22880
rect 15148 22816 15154 22880
rect 14838 22815 15154 22816
rect 21784 22880 22100 22881
rect 21784 22816 21790 22880
rect 21854 22816 21870 22880
rect 21934 22816 21950 22880
rect 22014 22816 22030 22880
rect 22094 22816 22100 22880
rect 21784 22815 22100 22816
rect 28730 22880 29046 22881
rect 28730 22816 28736 22880
rect 28800 22816 28816 22880
rect 28880 22816 28896 22880
rect 28960 22816 28976 22880
rect 29040 22816 29046 22880
rect 28730 22815 29046 22816
rect 4419 22336 4735 22337
rect 4419 22272 4425 22336
rect 4489 22272 4505 22336
rect 4569 22272 4585 22336
rect 4649 22272 4665 22336
rect 4729 22272 4735 22336
rect 4419 22271 4735 22272
rect 11365 22336 11681 22337
rect 11365 22272 11371 22336
rect 11435 22272 11451 22336
rect 11515 22272 11531 22336
rect 11595 22272 11611 22336
rect 11675 22272 11681 22336
rect 11365 22271 11681 22272
rect 18311 22336 18627 22337
rect 18311 22272 18317 22336
rect 18381 22272 18397 22336
rect 18461 22272 18477 22336
rect 18541 22272 18557 22336
rect 18621 22272 18627 22336
rect 18311 22271 18627 22272
rect 25257 22336 25573 22337
rect 25257 22272 25263 22336
rect 25327 22272 25343 22336
rect 25407 22272 25423 22336
rect 25487 22272 25503 22336
rect 25567 22272 25573 22336
rect 29200 22312 30000 22432
rect 25257 22271 25573 22272
rect 0 22130 800 22160
rect 1577 22130 1643 22133
rect 0 22128 1643 22130
rect 0 22072 1582 22128
rect 1638 22072 1643 22128
rect 0 22070 1643 22072
rect 0 22040 800 22070
rect 1577 22067 1643 22070
rect 28349 21994 28415 21997
rect 28349 21992 29378 21994
rect 28349 21936 28354 21992
rect 28410 21936 29378 21992
rect 28349 21934 29378 21936
rect 28349 21931 28415 21934
rect 7892 21792 8208 21793
rect 7892 21728 7898 21792
rect 7962 21728 7978 21792
rect 8042 21728 8058 21792
rect 8122 21728 8138 21792
rect 8202 21728 8208 21792
rect 7892 21727 8208 21728
rect 14838 21792 15154 21793
rect 14838 21728 14844 21792
rect 14908 21728 14924 21792
rect 14988 21728 15004 21792
rect 15068 21728 15084 21792
rect 15148 21728 15154 21792
rect 14838 21727 15154 21728
rect 21784 21792 22100 21793
rect 21784 21728 21790 21792
rect 21854 21728 21870 21792
rect 21934 21728 21950 21792
rect 22014 21728 22030 21792
rect 22094 21728 22100 21792
rect 21784 21727 22100 21728
rect 28730 21792 29046 21793
rect 28730 21728 28736 21792
rect 28800 21728 28816 21792
rect 28880 21728 28896 21792
rect 28960 21728 28976 21792
rect 29040 21728 29046 21792
rect 29318 21752 29378 21934
rect 28730 21727 29046 21728
rect 29200 21632 30000 21752
rect 0 21450 800 21480
rect 1577 21450 1643 21453
rect 0 21448 1643 21450
rect 0 21392 1582 21448
rect 1638 21392 1643 21448
rect 0 21390 1643 21392
rect 0 21360 800 21390
rect 1577 21387 1643 21390
rect 4419 21248 4735 21249
rect 4419 21184 4425 21248
rect 4489 21184 4505 21248
rect 4569 21184 4585 21248
rect 4649 21184 4665 21248
rect 4729 21184 4735 21248
rect 4419 21183 4735 21184
rect 11365 21248 11681 21249
rect 11365 21184 11371 21248
rect 11435 21184 11451 21248
rect 11515 21184 11531 21248
rect 11595 21184 11611 21248
rect 11675 21184 11681 21248
rect 11365 21183 11681 21184
rect 18311 21248 18627 21249
rect 18311 21184 18317 21248
rect 18381 21184 18397 21248
rect 18461 21184 18477 21248
rect 18541 21184 18557 21248
rect 18621 21184 18627 21248
rect 18311 21183 18627 21184
rect 25257 21248 25573 21249
rect 25257 21184 25263 21248
rect 25327 21184 25343 21248
rect 25407 21184 25423 21248
rect 25487 21184 25503 21248
rect 25567 21184 25573 21248
rect 25257 21183 25573 21184
rect 28349 21042 28415 21045
rect 29200 21042 30000 21072
rect 28349 21040 30000 21042
rect 28349 20984 28354 21040
rect 28410 20984 30000 21040
rect 28349 20982 30000 20984
rect 28349 20979 28415 20982
rect 29200 20952 30000 20982
rect 0 20680 800 20800
rect 7892 20704 8208 20705
rect 7892 20640 7898 20704
rect 7962 20640 7978 20704
rect 8042 20640 8058 20704
rect 8122 20640 8138 20704
rect 8202 20640 8208 20704
rect 7892 20639 8208 20640
rect 14838 20704 15154 20705
rect 14838 20640 14844 20704
rect 14908 20640 14924 20704
rect 14988 20640 15004 20704
rect 15068 20640 15084 20704
rect 15148 20640 15154 20704
rect 14838 20639 15154 20640
rect 21784 20704 22100 20705
rect 21784 20640 21790 20704
rect 21854 20640 21870 20704
rect 21934 20640 21950 20704
rect 22014 20640 22030 20704
rect 22094 20640 22100 20704
rect 21784 20639 22100 20640
rect 28730 20704 29046 20705
rect 28730 20640 28736 20704
rect 28800 20640 28816 20704
rect 28880 20640 28896 20704
rect 28960 20640 28976 20704
rect 29040 20640 29046 20704
rect 28730 20639 29046 20640
rect 29200 20272 30000 20392
rect 4419 20160 4735 20161
rect 0 20090 800 20120
rect 4419 20096 4425 20160
rect 4489 20096 4505 20160
rect 4569 20096 4585 20160
rect 4649 20096 4665 20160
rect 4729 20096 4735 20160
rect 4419 20095 4735 20096
rect 11365 20160 11681 20161
rect 11365 20096 11371 20160
rect 11435 20096 11451 20160
rect 11515 20096 11531 20160
rect 11595 20096 11611 20160
rect 11675 20096 11681 20160
rect 11365 20095 11681 20096
rect 18311 20160 18627 20161
rect 18311 20096 18317 20160
rect 18381 20096 18397 20160
rect 18461 20096 18477 20160
rect 18541 20096 18557 20160
rect 18621 20096 18627 20160
rect 18311 20095 18627 20096
rect 25257 20160 25573 20161
rect 25257 20096 25263 20160
rect 25327 20096 25343 20160
rect 25407 20096 25423 20160
rect 25487 20096 25503 20160
rect 25567 20096 25573 20160
rect 25257 20095 25573 20096
rect 1577 20090 1643 20093
rect 0 20088 1643 20090
rect 0 20032 1582 20088
rect 1638 20032 1643 20088
rect 0 20030 1643 20032
rect 0 20000 800 20030
rect 1577 20027 1643 20030
rect 28349 19954 28415 19957
rect 28349 19952 29378 19954
rect 28349 19896 28354 19952
rect 28410 19896 29378 19952
rect 28349 19894 29378 19896
rect 28349 19891 28415 19894
rect 29318 19712 29378 19894
rect 7892 19616 8208 19617
rect 7892 19552 7898 19616
rect 7962 19552 7978 19616
rect 8042 19552 8058 19616
rect 8122 19552 8138 19616
rect 8202 19552 8208 19616
rect 7892 19551 8208 19552
rect 14838 19616 15154 19617
rect 14838 19552 14844 19616
rect 14908 19552 14924 19616
rect 14988 19552 15004 19616
rect 15068 19552 15084 19616
rect 15148 19552 15154 19616
rect 14838 19551 15154 19552
rect 21784 19616 22100 19617
rect 21784 19552 21790 19616
rect 21854 19552 21870 19616
rect 21934 19552 21950 19616
rect 22014 19552 22030 19616
rect 22094 19552 22100 19616
rect 21784 19551 22100 19552
rect 28730 19616 29046 19617
rect 28730 19552 28736 19616
rect 28800 19552 28816 19616
rect 28880 19552 28896 19616
rect 28960 19552 28976 19616
rect 29040 19552 29046 19616
rect 29200 19592 30000 19712
rect 28730 19551 29046 19552
rect 0 19410 800 19440
rect 1577 19410 1643 19413
rect 0 19408 1643 19410
rect 0 19352 1582 19408
rect 1638 19352 1643 19408
rect 0 19350 1643 19352
rect 0 19320 800 19350
rect 1577 19347 1643 19350
rect 4419 19072 4735 19073
rect 4419 19008 4425 19072
rect 4489 19008 4505 19072
rect 4569 19008 4585 19072
rect 4649 19008 4665 19072
rect 4729 19008 4735 19072
rect 4419 19007 4735 19008
rect 11365 19072 11681 19073
rect 11365 19008 11371 19072
rect 11435 19008 11451 19072
rect 11515 19008 11531 19072
rect 11595 19008 11611 19072
rect 11675 19008 11681 19072
rect 11365 19007 11681 19008
rect 18311 19072 18627 19073
rect 18311 19008 18317 19072
rect 18381 19008 18397 19072
rect 18461 19008 18477 19072
rect 18541 19008 18557 19072
rect 18621 19008 18627 19072
rect 18311 19007 18627 19008
rect 25257 19072 25573 19073
rect 25257 19008 25263 19072
rect 25327 19008 25343 19072
rect 25407 19008 25423 19072
rect 25487 19008 25503 19072
rect 25567 19008 25573 19072
rect 25257 19007 25573 19008
rect 28349 19002 28415 19005
rect 29200 19002 30000 19032
rect 28349 19000 30000 19002
rect 28349 18944 28354 19000
rect 28410 18944 30000 19000
rect 28349 18942 30000 18944
rect 28349 18939 28415 18942
rect 29200 18912 30000 18942
rect 0 18640 800 18760
rect 7892 18528 8208 18529
rect 7892 18464 7898 18528
rect 7962 18464 7978 18528
rect 8042 18464 8058 18528
rect 8122 18464 8138 18528
rect 8202 18464 8208 18528
rect 7892 18463 8208 18464
rect 14838 18528 15154 18529
rect 14838 18464 14844 18528
rect 14908 18464 14924 18528
rect 14988 18464 15004 18528
rect 15068 18464 15084 18528
rect 15148 18464 15154 18528
rect 14838 18463 15154 18464
rect 21784 18528 22100 18529
rect 21784 18464 21790 18528
rect 21854 18464 21870 18528
rect 21934 18464 21950 18528
rect 22014 18464 22030 18528
rect 22094 18464 22100 18528
rect 21784 18463 22100 18464
rect 28730 18528 29046 18529
rect 28730 18464 28736 18528
rect 28800 18464 28816 18528
rect 28880 18464 28896 18528
rect 28960 18464 28976 18528
rect 29040 18464 29046 18528
rect 28730 18463 29046 18464
rect 29200 18232 30000 18352
rect 0 18050 800 18080
rect 1577 18050 1643 18053
rect 0 18048 1643 18050
rect 0 17992 1582 18048
rect 1638 17992 1643 18048
rect 0 17990 1643 17992
rect 0 17960 800 17990
rect 1577 17987 1643 17990
rect 4419 17984 4735 17985
rect 4419 17920 4425 17984
rect 4489 17920 4505 17984
rect 4569 17920 4585 17984
rect 4649 17920 4665 17984
rect 4729 17920 4735 17984
rect 4419 17919 4735 17920
rect 11365 17984 11681 17985
rect 11365 17920 11371 17984
rect 11435 17920 11451 17984
rect 11515 17920 11531 17984
rect 11595 17920 11611 17984
rect 11675 17920 11681 17984
rect 11365 17919 11681 17920
rect 18311 17984 18627 17985
rect 18311 17920 18317 17984
rect 18381 17920 18397 17984
rect 18461 17920 18477 17984
rect 18541 17920 18557 17984
rect 18621 17920 18627 17984
rect 18311 17919 18627 17920
rect 25257 17984 25573 17985
rect 25257 17920 25263 17984
rect 25327 17920 25343 17984
rect 25407 17920 25423 17984
rect 25487 17920 25503 17984
rect 25567 17920 25573 17984
rect 25257 17919 25573 17920
rect 28349 17642 28415 17645
rect 29200 17642 30000 17672
rect 28349 17640 30000 17642
rect 28349 17584 28354 17640
rect 28410 17584 30000 17640
rect 28349 17582 30000 17584
rect 28349 17579 28415 17582
rect 29200 17552 30000 17582
rect 7892 17440 8208 17441
rect 0 17370 800 17400
rect 7892 17376 7898 17440
rect 7962 17376 7978 17440
rect 8042 17376 8058 17440
rect 8122 17376 8138 17440
rect 8202 17376 8208 17440
rect 7892 17375 8208 17376
rect 14838 17440 15154 17441
rect 14838 17376 14844 17440
rect 14908 17376 14924 17440
rect 14988 17376 15004 17440
rect 15068 17376 15084 17440
rect 15148 17376 15154 17440
rect 14838 17375 15154 17376
rect 21784 17440 22100 17441
rect 21784 17376 21790 17440
rect 21854 17376 21870 17440
rect 21934 17376 21950 17440
rect 22014 17376 22030 17440
rect 22094 17376 22100 17440
rect 21784 17375 22100 17376
rect 28730 17440 29046 17441
rect 28730 17376 28736 17440
rect 28800 17376 28816 17440
rect 28880 17376 28896 17440
rect 28960 17376 28976 17440
rect 29040 17376 29046 17440
rect 28730 17375 29046 17376
rect 1577 17370 1643 17373
rect 0 17368 1643 17370
rect 0 17312 1582 17368
rect 1638 17312 1643 17368
rect 0 17310 1643 17312
rect 0 17280 800 17310
rect 1577 17307 1643 17310
rect 28349 16962 28415 16965
rect 29200 16962 30000 16992
rect 28349 16960 30000 16962
rect 28349 16904 28354 16960
rect 28410 16904 30000 16960
rect 28349 16902 30000 16904
rect 28349 16899 28415 16902
rect 4419 16896 4735 16897
rect 4419 16832 4425 16896
rect 4489 16832 4505 16896
rect 4569 16832 4585 16896
rect 4649 16832 4665 16896
rect 4729 16832 4735 16896
rect 4419 16831 4735 16832
rect 11365 16896 11681 16897
rect 11365 16832 11371 16896
rect 11435 16832 11451 16896
rect 11515 16832 11531 16896
rect 11595 16832 11611 16896
rect 11675 16832 11681 16896
rect 11365 16831 11681 16832
rect 18311 16896 18627 16897
rect 18311 16832 18317 16896
rect 18381 16832 18397 16896
rect 18461 16832 18477 16896
rect 18541 16832 18557 16896
rect 18621 16832 18627 16896
rect 18311 16831 18627 16832
rect 25257 16896 25573 16897
rect 25257 16832 25263 16896
rect 25327 16832 25343 16896
rect 25407 16832 25423 16896
rect 25487 16832 25503 16896
rect 25567 16832 25573 16896
rect 29200 16872 30000 16902
rect 25257 16831 25573 16832
rect 0 16600 800 16720
rect 7892 16352 8208 16353
rect 7892 16288 7898 16352
rect 7962 16288 7978 16352
rect 8042 16288 8058 16352
rect 8122 16288 8138 16352
rect 8202 16288 8208 16352
rect 7892 16287 8208 16288
rect 14838 16352 15154 16353
rect 14838 16288 14844 16352
rect 14908 16288 14924 16352
rect 14988 16288 15004 16352
rect 15068 16288 15084 16352
rect 15148 16288 15154 16352
rect 14838 16287 15154 16288
rect 21784 16352 22100 16353
rect 21784 16288 21790 16352
rect 21854 16288 21870 16352
rect 21934 16288 21950 16352
rect 22014 16288 22030 16352
rect 22094 16288 22100 16352
rect 21784 16287 22100 16288
rect 28730 16352 29046 16353
rect 28730 16288 28736 16352
rect 28800 16288 28816 16352
rect 28880 16288 28896 16352
rect 28960 16288 28976 16352
rect 29040 16288 29046 16352
rect 28730 16287 29046 16288
rect 29200 16192 30000 16312
rect 0 16010 800 16040
rect 1577 16010 1643 16013
rect 0 16008 1643 16010
rect 0 15952 1582 16008
rect 1638 15952 1643 16008
rect 0 15950 1643 15952
rect 0 15920 800 15950
rect 1577 15947 1643 15950
rect 4419 15808 4735 15809
rect 4419 15744 4425 15808
rect 4489 15744 4505 15808
rect 4569 15744 4585 15808
rect 4649 15744 4665 15808
rect 4729 15744 4735 15808
rect 4419 15743 4735 15744
rect 11365 15808 11681 15809
rect 11365 15744 11371 15808
rect 11435 15744 11451 15808
rect 11515 15744 11531 15808
rect 11595 15744 11611 15808
rect 11675 15744 11681 15808
rect 11365 15743 11681 15744
rect 18311 15808 18627 15809
rect 18311 15744 18317 15808
rect 18381 15744 18397 15808
rect 18461 15744 18477 15808
rect 18541 15744 18557 15808
rect 18621 15744 18627 15808
rect 18311 15743 18627 15744
rect 25257 15808 25573 15809
rect 25257 15744 25263 15808
rect 25327 15744 25343 15808
rect 25407 15744 25423 15808
rect 25487 15744 25503 15808
rect 25567 15744 25573 15808
rect 25257 15743 25573 15744
rect 28349 15602 28415 15605
rect 29200 15602 30000 15632
rect 28349 15600 30000 15602
rect 28349 15544 28354 15600
rect 28410 15544 30000 15600
rect 28349 15542 30000 15544
rect 28349 15539 28415 15542
rect 29200 15512 30000 15542
rect 0 15330 800 15360
rect 1577 15330 1643 15333
rect 0 15328 1643 15330
rect 0 15272 1582 15328
rect 1638 15272 1643 15328
rect 0 15270 1643 15272
rect 0 15240 800 15270
rect 1577 15267 1643 15270
rect 7892 15264 8208 15265
rect 7892 15200 7898 15264
rect 7962 15200 7978 15264
rect 8042 15200 8058 15264
rect 8122 15200 8138 15264
rect 8202 15200 8208 15264
rect 7892 15199 8208 15200
rect 14838 15264 15154 15265
rect 14838 15200 14844 15264
rect 14908 15200 14924 15264
rect 14988 15200 15004 15264
rect 15068 15200 15084 15264
rect 15148 15200 15154 15264
rect 14838 15199 15154 15200
rect 21784 15264 22100 15265
rect 21784 15200 21790 15264
rect 21854 15200 21870 15264
rect 21934 15200 21950 15264
rect 22014 15200 22030 15264
rect 22094 15200 22100 15264
rect 21784 15199 22100 15200
rect 28730 15264 29046 15265
rect 28730 15200 28736 15264
rect 28800 15200 28816 15264
rect 28880 15200 28896 15264
rect 28960 15200 28976 15264
rect 29040 15200 29046 15264
rect 28730 15199 29046 15200
rect 28349 14922 28415 14925
rect 29200 14922 30000 14952
rect 28349 14920 30000 14922
rect 28349 14864 28354 14920
rect 28410 14864 30000 14920
rect 28349 14862 30000 14864
rect 28349 14859 28415 14862
rect 29200 14832 30000 14862
rect 4419 14720 4735 14721
rect 0 14560 800 14680
rect 4419 14656 4425 14720
rect 4489 14656 4505 14720
rect 4569 14656 4585 14720
rect 4649 14656 4665 14720
rect 4729 14656 4735 14720
rect 4419 14655 4735 14656
rect 11365 14720 11681 14721
rect 11365 14656 11371 14720
rect 11435 14656 11451 14720
rect 11515 14656 11531 14720
rect 11595 14656 11611 14720
rect 11675 14656 11681 14720
rect 11365 14655 11681 14656
rect 18311 14720 18627 14721
rect 18311 14656 18317 14720
rect 18381 14656 18397 14720
rect 18461 14656 18477 14720
rect 18541 14656 18557 14720
rect 18621 14656 18627 14720
rect 18311 14655 18627 14656
rect 25257 14720 25573 14721
rect 25257 14656 25263 14720
rect 25327 14656 25343 14720
rect 25407 14656 25423 14720
rect 25487 14656 25503 14720
rect 25567 14656 25573 14720
rect 25257 14655 25573 14656
rect 7892 14176 8208 14177
rect 7892 14112 7898 14176
rect 7962 14112 7978 14176
rect 8042 14112 8058 14176
rect 8122 14112 8138 14176
rect 8202 14112 8208 14176
rect 7892 14111 8208 14112
rect 14838 14176 15154 14177
rect 14838 14112 14844 14176
rect 14908 14112 14924 14176
rect 14988 14112 15004 14176
rect 15068 14112 15084 14176
rect 15148 14112 15154 14176
rect 14838 14111 15154 14112
rect 21784 14176 22100 14177
rect 21784 14112 21790 14176
rect 21854 14112 21870 14176
rect 21934 14112 21950 14176
rect 22014 14112 22030 14176
rect 22094 14112 22100 14176
rect 21784 14111 22100 14112
rect 28730 14176 29046 14177
rect 28730 14112 28736 14176
rect 28800 14112 28816 14176
rect 28880 14112 28896 14176
rect 28960 14112 28976 14176
rect 29040 14112 29046 14176
rect 29200 14152 30000 14272
rect 28730 14111 29046 14112
rect 0 13970 800 14000
rect 1577 13970 1643 13973
rect 0 13968 1643 13970
rect 0 13912 1582 13968
rect 1638 13912 1643 13968
rect 0 13910 1643 13912
rect 0 13880 800 13910
rect 1577 13907 1643 13910
rect 4419 13632 4735 13633
rect 4419 13568 4425 13632
rect 4489 13568 4505 13632
rect 4569 13568 4585 13632
rect 4649 13568 4665 13632
rect 4729 13568 4735 13632
rect 4419 13567 4735 13568
rect 11365 13632 11681 13633
rect 11365 13568 11371 13632
rect 11435 13568 11451 13632
rect 11515 13568 11531 13632
rect 11595 13568 11611 13632
rect 11675 13568 11681 13632
rect 11365 13567 11681 13568
rect 18311 13632 18627 13633
rect 18311 13568 18317 13632
rect 18381 13568 18397 13632
rect 18461 13568 18477 13632
rect 18541 13568 18557 13632
rect 18621 13568 18627 13632
rect 18311 13567 18627 13568
rect 25257 13632 25573 13633
rect 25257 13568 25263 13632
rect 25327 13568 25343 13632
rect 25407 13568 25423 13632
rect 25487 13568 25503 13632
rect 25567 13568 25573 13632
rect 25257 13567 25573 13568
rect 28349 13562 28415 13565
rect 29200 13562 30000 13592
rect 28349 13560 30000 13562
rect 28349 13504 28354 13560
rect 28410 13504 30000 13560
rect 28349 13502 30000 13504
rect 28349 13499 28415 13502
rect 29200 13472 30000 13502
rect 0 13290 800 13320
rect 1577 13290 1643 13293
rect 0 13288 1643 13290
rect 0 13232 1582 13288
rect 1638 13232 1643 13288
rect 0 13230 1643 13232
rect 0 13200 800 13230
rect 1577 13227 1643 13230
rect 7892 13088 8208 13089
rect 7892 13024 7898 13088
rect 7962 13024 7978 13088
rect 8042 13024 8058 13088
rect 8122 13024 8138 13088
rect 8202 13024 8208 13088
rect 7892 13023 8208 13024
rect 14838 13088 15154 13089
rect 14838 13024 14844 13088
rect 14908 13024 14924 13088
rect 14988 13024 15004 13088
rect 15068 13024 15084 13088
rect 15148 13024 15154 13088
rect 14838 13023 15154 13024
rect 21784 13088 22100 13089
rect 21784 13024 21790 13088
rect 21854 13024 21870 13088
rect 21934 13024 21950 13088
rect 22014 13024 22030 13088
rect 22094 13024 22100 13088
rect 21784 13023 22100 13024
rect 28730 13088 29046 13089
rect 28730 13024 28736 13088
rect 28800 13024 28816 13088
rect 28880 13024 28896 13088
rect 28960 13024 28976 13088
rect 29040 13024 29046 13088
rect 28730 13023 29046 13024
rect 28349 12882 28415 12885
rect 29200 12882 30000 12912
rect 28349 12880 30000 12882
rect 28349 12824 28354 12880
rect 28410 12824 30000 12880
rect 28349 12822 30000 12824
rect 28349 12819 28415 12822
rect 29200 12792 30000 12822
rect 0 12520 800 12640
rect 4419 12544 4735 12545
rect 4419 12480 4425 12544
rect 4489 12480 4505 12544
rect 4569 12480 4585 12544
rect 4649 12480 4665 12544
rect 4729 12480 4735 12544
rect 4419 12479 4735 12480
rect 11365 12544 11681 12545
rect 11365 12480 11371 12544
rect 11435 12480 11451 12544
rect 11515 12480 11531 12544
rect 11595 12480 11611 12544
rect 11675 12480 11681 12544
rect 11365 12479 11681 12480
rect 18311 12544 18627 12545
rect 18311 12480 18317 12544
rect 18381 12480 18397 12544
rect 18461 12480 18477 12544
rect 18541 12480 18557 12544
rect 18621 12480 18627 12544
rect 18311 12479 18627 12480
rect 25257 12544 25573 12545
rect 25257 12480 25263 12544
rect 25327 12480 25343 12544
rect 25407 12480 25423 12544
rect 25487 12480 25503 12544
rect 25567 12480 25573 12544
rect 25257 12479 25573 12480
rect 29200 12112 30000 12232
rect 7892 12000 8208 12001
rect 0 11930 800 11960
rect 7892 11936 7898 12000
rect 7962 11936 7978 12000
rect 8042 11936 8058 12000
rect 8122 11936 8138 12000
rect 8202 11936 8208 12000
rect 7892 11935 8208 11936
rect 14838 12000 15154 12001
rect 14838 11936 14844 12000
rect 14908 11936 14924 12000
rect 14988 11936 15004 12000
rect 15068 11936 15084 12000
rect 15148 11936 15154 12000
rect 14838 11935 15154 11936
rect 21784 12000 22100 12001
rect 21784 11936 21790 12000
rect 21854 11936 21870 12000
rect 21934 11936 21950 12000
rect 22014 11936 22030 12000
rect 22094 11936 22100 12000
rect 21784 11935 22100 11936
rect 28730 12000 29046 12001
rect 28730 11936 28736 12000
rect 28800 11936 28816 12000
rect 28880 11936 28896 12000
rect 28960 11936 28976 12000
rect 29040 11936 29046 12000
rect 28730 11935 29046 11936
rect 1577 11930 1643 11933
rect 0 11928 1643 11930
rect 0 11872 1582 11928
rect 1638 11872 1643 11928
rect 0 11870 1643 11872
rect 0 11840 800 11870
rect 1577 11867 1643 11870
rect 28349 11522 28415 11525
rect 29200 11522 30000 11552
rect 28349 11520 30000 11522
rect 28349 11464 28354 11520
rect 28410 11464 30000 11520
rect 28349 11462 30000 11464
rect 28349 11459 28415 11462
rect 4419 11456 4735 11457
rect 4419 11392 4425 11456
rect 4489 11392 4505 11456
rect 4569 11392 4585 11456
rect 4649 11392 4665 11456
rect 4729 11392 4735 11456
rect 4419 11391 4735 11392
rect 11365 11456 11681 11457
rect 11365 11392 11371 11456
rect 11435 11392 11451 11456
rect 11515 11392 11531 11456
rect 11595 11392 11611 11456
rect 11675 11392 11681 11456
rect 11365 11391 11681 11392
rect 18311 11456 18627 11457
rect 18311 11392 18317 11456
rect 18381 11392 18397 11456
rect 18461 11392 18477 11456
rect 18541 11392 18557 11456
rect 18621 11392 18627 11456
rect 18311 11391 18627 11392
rect 25257 11456 25573 11457
rect 25257 11392 25263 11456
rect 25327 11392 25343 11456
rect 25407 11392 25423 11456
rect 25487 11392 25503 11456
rect 25567 11392 25573 11456
rect 29200 11432 30000 11462
rect 25257 11391 25573 11392
rect 0 11250 800 11280
rect 1577 11250 1643 11253
rect 0 11248 1643 11250
rect 0 11192 1582 11248
rect 1638 11192 1643 11248
rect 0 11190 1643 11192
rect 0 11160 800 11190
rect 1577 11187 1643 11190
rect 28349 11114 28415 11117
rect 28349 11112 29378 11114
rect 28349 11056 28354 11112
rect 28410 11056 29378 11112
rect 28349 11054 29378 11056
rect 28349 11051 28415 11054
rect 7892 10912 8208 10913
rect 7892 10848 7898 10912
rect 7962 10848 7978 10912
rect 8042 10848 8058 10912
rect 8122 10848 8138 10912
rect 8202 10848 8208 10912
rect 7892 10847 8208 10848
rect 14838 10912 15154 10913
rect 14838 10848 14844 10912
rect 14908 10848 14924 10912
rect 14988 10848 15004 10912
rect 15068 10848 15084 10912
rect 15148 10848 15154 10912
rect 14838 10847 15154 10848
rect 21784 10912 22100 10913
rect 21784 10848 21790 10912
rect 21854 10848 21870 10912
rect 21934 10848 21950 10912
rect 22014 10848 22030 10912
rect 22094 10848 22100 10912
rect 21784 10847 22100 10848
rect 28730 10912 29046 10913
rect 28730 10848 28736 10912
rect 28800 10848 28816 10912
rect 28880 10848 28896 10912
rect 28960 10848 28976 10912
rect 29040 10848 29046 10912
rect 29318 10872 29378 11054
rect 28730 10847 29046 10848
rect 29200 10752 30000 10872
rect 0 10480 800 10600
rect 4419 10368 4735 10369
rect 4419 10304 4425 10368
rect 4489 10304 4505 10368
rect 4569 10304 4585 10368
rect 4649 10304 4665 10368
rect 4729 10304 4735 10368
rect 4419 10303 4735 10304
rect 11365 10368 11681 10369
rect 11365 10304 11371 10368
rect 11435 10304 11451 10368
rect 11515 10304 11531 10368
rect 11595 10304 11611 10368
rect 11675 10304 11681 10368
rect 11365 10303 11681 10304
rect 18311 10368 18627 10369
rect 18311 10304 18317 10368
rect 18381 10304 18397 10368
rect 18461 10304 18477 10368
rect 18541 10304 18557 10368
rect 18621 10304 18627 10368
rect 18311 10303 18627 10304
rect 25257 10368 25573 10369
rect 25257 10304 25263 10368
rect 25327 10304 25343 10368
rect 25407 10304 25423 10368
rect 25487 10304 25503 10368
rect 25567 10304 25573 10368
rect 25257 10303 25573 10304
rect 29200 10072 30000 10192
rect 0 9890 800 9920
rect 1577 9890 1643 9893
rect 0 9888 1643 9890
rect 0 9832 1582 9888
rect 1638 9832 1643 9888
rect 0 9830 1643 9832
rect 0 9800 800 9830
rect 1577 9827 1643 9830
rect 7892 9824 8208 9825
rect 7892 9760 7898 9824
rect 7962 9760 7978 9824
rect 8042 9760 8058 9824
rect 8122 9760 8138 9824
rect 8202 9760 8208 9824
rect 7892 9759 8208 9760
rect 14838 9824 15154 9825
rect 14838 9760 14844 9824
rect 14908 9760 14924 9824
rect 14988 9760 15004 9824
rect 15068 9760 15084 9824
rect 15148 9760 15154 9824
rect 14838 9759 15154 9760
rect 21784 9824 22100 9825
rect 21784 9760 21790 9824
rect 21854 9760 21870 9824
rect 21934 9760 21950 9824
rect 22014 9760 22030 9824
rect 22094 9760 22100 9824
rect 21784 9759 22100 9760
rect 28730 9824 29046 9825
rect 28730 9760 28736 9824
rect 28800 9760 28816 9824
rect 28880 9760 28896 9824
rect 28960 9760 28976 9824
rect 29040 9760 29046 9824
rect 28730 9759 29046 9760
rect 28349 9482 28415 9485
rect 29200 9482 30000 9512
rect 28349 9480 30000 9482
rect 28349 9424 28354 9480
rect 28410 9424 30000 9480
rect 28349 9422 30000 9424
rect 28349 9419 28415 9422
rect 29200 9392 30000 9422
rect 4419 9280 4735 9281
rect 0 9210 800 9240
rect 4419 9216 4425 9280
rect 4489 9216 4505 9280
rect 4569 9216 4585 9280
rect 4649 9216 4665 9280
rect 4729 9216 4735 9280
rect 4419 9215 4735 9216
rect 11365 9280 11681 9281
rect 11365 9216 11371 9280
rect 11435 9216 11451 9280
rect 11515 9216 11531 9280
rect 11595 9216 11611 9280
rect 11675 9216 11681 9280
rect 11365 9215 11681 9216
rect 18311 9280 18627 9281
rect 18311 9216 18317 9280
rect 18381 9216 18397 9280
rect 18461 9216 18477 9280
rect 18541 9216 18557 9280
rect 18621 9216 18627 9280
rect 18311 9215 18627 9216
rect 25257 9280 25573 9281
rect 25257 9216 25263 9280
rect 25327 9216 25343 9280
rect 25407 9216 25423 9280
rect 25487 9216 25503 9280
rect 25567 9216 25573 9280
rect 25257 9215 25573 9216
rect 1577 9210 1643 9213
rect 0 9208 1643 9210
rect 0 9152 1582 9208
rect 1638 9152 1643 9208
rect 0 9150 1643 9152
rect 0 9120 800 9150
rect 1577 9147 1643 9150
rect 28349 9074 28415 9077
rect 28349 9072 29378 9074
rect 28349 9016 28354 9072
rect 28410 9016 29378 9072
rect 28349 9014 29378 9016
rect 28349 9011 28415 9014
rect 29318 8832 29378 9014
rect 7892 8736 8208 8737
rect 7892 8672 7898 8736
rect 7962 8672 7978 8736
rect 8042 8672 8058 8736
rect 8122 8672 8138 8736
rect 8202 8672 8208 8736
rect 7892 8671 8208 8672
rect 14838 8736 15154 8737
rect 14838 8672 14844 8736
rect 14908 8672 14924 8736
rect 14988 8672 15004 8736
rect 15068 8672 15084 8736
rect 15148 8672 15154 8736
rect 14838 8671 15154 8672
rect 21784 8736 22100 8737
rect 21784 8672 21790 8736
rect 21854 8672 21870 8736
rect 21934 8672 21950 8736
rect 22014 8672 22030 8736
rect 22094 8672 22100 8736
rect 21784 8671 22100 8672
rect 28730 8736 29046 8737
rect 28730 8672 28736 8736
rect 28800 8672 28816 8736
rect 28880 8672 28896 8736
rect 28960 8672 28976 8736
rect 29040 8672 29046 8736
rect 29200 8712 30000 8832
rect 28730 8671 29046 8672
rect 0 8440 800 8560
rect 4419 8192 4735 8193
rect 4419 8128 4425 8192
rect 4489 8128 4505 8192
rect 4569 8128 4585 8192
rect 4649 8128 4665 8192
rect 4729 8128 4735 8192
rect 4419 8127 4735 8128
rect 11365 8192 11681 8193
rect 11365 8128 11371 8192
rect 11435 8128 11451 8192
rect 11515 8128 11531 8192
rect 11595 8128 11611 8192
rect 11675 8128 11681 8192
rect 11365 8127 11681 8128
rect 18311 8192 18627 8193
rect 18311 8128 18317 8192
rect 18381 8128 18397 8192
rect 18461 8128 18477 8192
rect 18541 8128 18557 8192
rect 18621 8128 18627 8192
rect 18311 8127 18627 8128
rect 25257 8192 25573 8193
rect 25257 8128 25263 8192
rect 25327 8128 25343 8192
rect 25407 8128 25423 8192
rect 25487 8128 25503 8192
rect 25567 8128 25573 8192
rect 25257 8127 25573 8128
rect 29200 8032 30000 8152
rect 0 7850 800 7880
rect 1577 7850 1643 7853
rect 0 7848 1643 7850
rect 0 7792 1582 7848
rect 1638 7792 1643 7848
rect 0 7790 1643 7792
rect 0 7760 800 7790
rect 1577 7787 1643 7790
rect 7892 7648 8208 7649
rect 7892 7584 7898 7648
rect 7962 7584 7978 7648
rect 8042 7584 8058 7648
rect 8122 7584 8138 7648
rect 8202 7584 8208 7648
rect 7892 7583 8208 7584
rect 14838 7648 15154 7649
rect 14838 7584 14844 7648
rect 14908 7584 14924 7648
rect 14988 7584 15004 7648
rect 15068 7584 15084 7648
rect 15148 7584 15154 7648
rect 14838 7583 15154 7584
rect 21784 7648 22100 7649
rect 21784 7584 21790 7648
rect 21854 7584 21870 7648
rect 21934 7584 21950 7648
rect 22014 7584 22030 7648
rect 22094 7584 22100 7648
rect 21784 7583 22100 7584
rect 28730 7648 29046 7649
rect 28730 7584 28736 7648
rect 28800 7584 28816 7648
rect 28880 7584 28896 7648
rect 28960 7584 28976 7648
rect 29040 7584 29046 7648
rect 28730 7583 29046 7584
rect 28349 7442 28415 7445
rect 29200 7442 30000 7472
rect 28349 7440 30000 7442
rect 28349 7384 28354 7440
rect 28410 7384 30000 7440
rect 28349 7382 30000 7384
rect 28349 7379 28415 7382
rect 29200 7352 30000 7382
rect 0 7170 800 7200
rect 1577 7170 1643 7173
rect 0 7168 1643 7170
rect 0 7112 1582 7168
rect 1638 7112 1643 7168
rect 0 7110 1643 7112
rect 0 7080 800 7110
rect 1577 7107 1643 7110
rect 4419 7104 4735 7105
rect 4419 7040 4425 7104
rect 4489 7040 4505 7104
rect 4569 7040 4585 7104
rect 4649 7040 4665 7104
rect 4729 7040 4735 7104
rect 4419 7039 4735 7040
rect 11365 7104 11681 7105
rect 11365 7040 11371 7104
rect 11435 7040 11451 7104
rect 11515 7040 11531 7104
rect 11595 7040 11611 7104
rect 11675 7040 11681 7104
rect 11365 7039 11681 7040
rect 18311 7104 18627 7105
rect 18311 7040 18317 7104
rect 18381 7040 18397 7104
rect 18461 7040 18477 7104
rect 18541 7040 18557 7104
rect 18621 7040 18627 7104
rect 18311 7039 18627 7040
rect 25257 7104 25573 7105
rect 25257 7040 25263 7104
rect 25327 7040 25343 7104
rect 25407 7040 25423 7104
rect 25487 7040 25503 7104
rect 25567 7040 25573 7104
rect 25257 7039 25573 7040
rect 28349 6762 28415 6765
rect 29200 6762 30000 6792
rect 28349 6760 30000 6762
rect 28349 6704 28354 6760
rect 28410 6704 30000 6760
rect 28349 6702 30000 6704
rect 28349 6699 28415 6702
rect 29200 6672 30000 6702
rect 7892 6560 8208 6561
rect 0 6400 800 6520
rect 7892 6496 7898 6560
rect 7962 6496 7978 6560
rect 8042 6496 8058 6560
rect 8122 6496 8138 6560
rect 8202 6496 8208 6560
rect 7892 6495 8208 6496
rect 14838 6560 15154 6561
rect 14838 6496 14844 6560
rect 14908 6496 14924 6560
rect 14988 6496 15004 6560
rect 15068 6496 15084 6560
rect 15148 6496 15154 6560
rect 14838 6495 15154 6496
rect 21784 6560 22100 6561
rect 21784 6496 21790 6560
rect 21854 6496 21870 6560
rect 21934 6496 21950 6560
rect 22014 6496 22030 6560
rect 22094 6496 22100 6560
rect 21784 6495 22100 6496
rect 28730 6560 29046 6561
rect 28730 6496 28736 6560
rect 28800 6496 28816 6560
rect 28880 6496 28896 6560
rect 28960 6496 28976 6560
rect 29040 6496 29046 6560
rect 28730 6495 29046 6496
rect 4419 6016 4735 6017
rect 4419 5952 4425 6016
rect 4489 5952 4505 6016
rect 4569 5952 4585 6016
rect 4649 5952 4665 6016
rect 4729 5952 4735 6016
rect 4419 5951 4735 5952
rect 11365 6016 11681 6017
rect 11365 5952 11371 6016
rect 11435 5952 11451 6016
rect 11515 5952 11531 6016
rect 11595 5952 11611 6016
rect 11675 5952 11681 6016
rect 11365 5951 11681 5952
rect 18311 6016 18627 6017
rect 18311 5952 18317 6016
rect 18381 5952 18397 6016
rect 18461 5952 18477 6016
rect 18541 5952 18557 6016
rect 18621 5952 18627 6016
rect 18311 5951 18627 5952
rect 25257 6016 25573 6017
rect 25257 5952 25263 6016
rect 25327 5952 25343 6016
rect 25407 5952 25423 6016
rect 25487 5952 25503 6016
rect 25567 5952 25573 6016
rect 29200 5992 30000 6112
rect 25257 5951 25573 5952
rect 0 5810 800 5840
rect 1577 5810 1643 5813
rect 0 5808 1643 5810
rect 0 5752 1582 5808
rect 1638 5752 1643 5808
rect 0 5750 1643 5752
rect 0 5720 800 5750
rect 1577 5747 1643 5750
rect 28349 5674 28415 5677
rect 28349 5672 29378 5674
rect 28349 5616 28354 5672
rect 28410 5616 29378 5672
rect 28349 5614 29378 5616
rect 28349 5611 28415 5614
rect 7892 5472 8208 5473
rect 7892 5408 7898 5472
rect 7962 5408 7978 5472
rect 8042 5408 8058 5472
rect 8122 5408 8138 5472
rect 8202 5408 8208 5472
rect 7892 5407 8208 5408
rect 14838 5472 15154 5473
rect 14838 5408 14844 5472
rect 14908 5408 14924 5472
rect 14988 5408 15004 5472
rect 15068 5408 15084 5472
rect 15148 5408 15154 5472
rect 14838 5407 15154 5408
rect 21784 5472 22100 5473
rect 21784 5408 21790 5472
rect 21854 5408 21870 5472
rect 21934 5408 21950 5472
rect 22014 5408 22030 5472
rect 22094 5408 22100 5472
rect 21784 5407 22100 5408
rect 28730 5472 29046 5473
rect 28730 5408 28736 5472
rect 28800 5408 28816 5472
rect 28880 5408 28896 5472
rect 28960 5408 28976 5472
rect 29040 5408 29046 5472
rect 29318 5432 29378 5614
rect 28730 5407 29046 5408
rect 29200 5312 30000 5432
rect 0 5130 800 5160
rect 1577 5130 1643 5133
rect 0 5128 1643 5130
rect 0 5072 1582 5128
rect 1638 5072 1643 5128
rect 0 5070 1643 5072
rect 0 5040 800 5070
rect 1577 5067 1643 5070
rect 4419 4928 4735 4929
rect 4419 4864 4425 4928
rect 4489 4864 4505 4928
rect 4569 4864 4585 4928
rect 4649 4864 4665 4928
rect 4729 4864 4735 4928
rect 4419 4863 4735 4864
rect 11365 4928 11681 4929
rect 11365 4864 11371 4928
rect 11435 4864 11451 4928
rect 11515 4864 11531 4928
rect 11595 4864 11611 4928
rect 11675 4864 11681 4928
rect 11365 4863 11681 4864
rect 18311 4928 18627 4929
rect 18311 4864 18317 4928
rect 18381 4864 18397 4928
rect 18461 4864 18477 4928
rect 18541 4864 18557 4928
rect 18621 4864 18627 4928
rect 18311 4863 18627 4864
rect 25257 4928 25573 4929
rect 25257 4864 25263 4928
rect 25327 4864 25343 4928
rect 25407 4864 25423 4928
rect 25487 4864 25503 4928
rect 25567 4864 25573 4928
rect 25257 4863 25573 4864
rect 28349 4722 28415 4725
rect 29200 4722 30000 4752
rect 28349 4720 30000 4722
rect 28349 4664 28354 4720
rect 28410 4664 30000 4720
rect 28349 4662 30000 4664
rect 28349 4659 28415 4662
rect 29200 4632 30000 4662
rect 0 4360 800 4480
rect 7892 4384 8208 4385
rect 7892 4320 7898 4384
rect 7962 4320 7978 4384
rect 8042 4320 8058 4384
rect 8122 4320 8138 4384
rect 8202 4320 8208 4384
rect 7892 4319 8208 4320
rect 14838 4384 15154 4385
rect 14838 4320 14844 4384
rect 14908 4320 14924 4384
rect 14988 4320 15004 4384
rect 15068 4320 15084 4384
rect 15148 4320 15154 4384
rect 14838 4319 15154 4320
rect 21784 4384 22100 4385
rect 21784 4320 21790 4384
rect 21854 4320 21870 4384
rect 21934 4320 21950 4384
rect 22014 4320 22030 4384
rect 22094 4320 22100 4384
rect 21784 4319 22100 4320
rect 28730 4384 29046 4385
rect 28730 4320 28736 4384
rect 28800 4320 28816 4384
rect 28880 4320 28896 4384
rect 28960 4320 28976 4384
rect 29040 4320 29046 4384
rect 28730 4319 29046 4320
rect 28349 4042 28415 4045
rect 29200 4042 30000 4072
rect 28349 4040 30000 4042
rect 28349 3984 28354 4040
rect 28410 3984 30000 4040
rect 28349 3982 30000 3984
rect 28349 3979 28415 3982
rect 29200 3952 30000 3982
rect 4419 3840 4735 3841
rect 0 3770 800 3800
rect 4419 3776 4425 3840
rect 4489 3776 4505 3840
rect 4569 3776 4585 3840
rect 4649 3776 4665 3840
rect 4729 3776 4735 3840
rect 4419 3775 4735 3776
rect 11365 3840 11681 3841
rect 11365 3776 11371 3840
rect 11435 3776 11451 3840
rect 11515 3776 11531 3840
rect 11595 3776 11611 3840
rect 11675 3776 11681 3840
rect 11365 3775 11681 3776
rect 18311 3840 18627 3841
rect 18311 3776 18317 3840
rect 18381 3776 18397 3840
rect 18461 3776 18477 3840
rect 18541 3776 18557 3840
rect 18621 3776 18627 3840
rect 18311 3775 18627 3776
rect 25257 3840 25573 3841
rect 25257 3776 25263 3840
rect 25327 3776 25343 3840
rect 25407 3776 25423 3840
rect 25487 3776 25503 3840
rect 25567 3776 25573 3840
rect 25257 3775 25573 3776
rect 1577 3770 1643 3773
rect 0 3768 1643 3770
rect 0 3712 1582 3768
rect 1638 3712 1643 3768
rect 0 3710 1643 3712
rect 0 3680 800 3710
rect 1577 3707 1643 3710
rect 28349 3634 28415 3637
rect 28349 3632 29378 3634
rect 28349 3576 28354 3632
rect 28410 3576 29378 3632
rect 28349 3574 29378 3576
rect 28349 3571 28415 3574
rect 29318 3392 29378 3574
rect 7892 3296 8208 3297
rect 7892 3232 7898 3296
rect 7962 3232 7978 3296
rect 8042 3232 8058 3296
rect 8122 3232 8138 3296
rect 8202 3232 8208 3296
rect 7892 3231 8208 3232
rect 14838 3296 15154 3297
rect 14838 3232 14844 3296
rect 14908 3232 14924 3296
rect 14988 3232 15004 3296
rect 15068 3232 15084 3296
rect 15148 3232 15154 3296
rect 14838 3231 15154 3232
rect 21784 3296 22100 3297
rect 21784 3232 21790 3296
rect 21854 3232 21870 3296
rect 21934 3232 21950 3296
rect 22014 3232 22030 3296
rect 22094 3232 22100 3296
rect 21784 3231 22100 3232
rect 28730 3296 29046 3297
rect 28730 3232 28736 3296
rect 28800 3232 28816 3296
rect 28880 3232 28896 3296
rect 28960 3232 28976 3296
rect 29040 3232 29046 3296
rect 29200 3272 30000 3392
rect 28730 3231 29046 3232
rect 0 3090 800 3120
rect 1577 3090 1643 3093
rect 0 3088 1643 3090
rect 0 3032 1582 3088
rect 1638 3032 1643 3088
rect 0 3030 1643 3032
rect 0 3000 800 3030
rect 1577 3027 1643 3030
rect 4419 2752 4735 2753
rect 4419 2688 4425 2752
rect 4489 2688 4505 2752
rect 4569 2688 4585 2752
rect 4649 2688 4665 2752
rect 4729 2688 4735 2752
rect 4419 2687 4735 2688
rect 11365 2752 11681 2753
rect 11365 2688 11371 2752
rect 11435 2688 11451 2752
rect 11515 2688 11531 2752
rect 11595 2688 11611 2752
rect 11675 2688 11681 2752
rect 11365 2687 11681 2688
rect 18311 2752 18627 2753
rect 18311 2688 18317 2752
rect 18381 2688 18397 2752
rect 18461 2688 18477 2752
rect 18541 2688 18557 2752
rect 18621 2688 18627 2752
rect 18311 2687 18627 2688
rect 25257 2752 25573 2753
rect 25257 2688 25263 2752
rect 25327 2688 25343 2752
rect 25407 2688 25423 2752
rect 25487 2688 25503 2752
rect 25567 2688 25573 2752
rect 25257 2687 25573 2688
rect 28349 2682 28415 2685
rect 29200 2682 30000 2712
rect 28349 2680 30000 2682
rect 28349 2624 28354 2680
rect 28410 2624 30000 2680
rect 28349 2622 30000 2624
rect 28349 2619 28415 2622
rect 29200 2592 30000 2622
rect 7892 2208 8208 2209
rect 7892 2144 7898 2208
rect 7962 2144 7978 2208
rect 8042 2144 8058 2208
rect 8122 2144 8138 2208
rect 8202 2144 8208 2208
rect 7892 2143 8208 2144
rect 14838 2208 15154 2209
rect 14838 2144 14844 2208
rect 14908 2144 14924 2208
rect 14988 2144 15004 2208
rect 15068 2144 15084 2208
rect 15148 2144 15154 2208
rect 14838 2143 15154 2144
rect 21784 2208 22100 2209
rect 21784 2144 21790 2208
rect 21854 2144 21870 2208
rect 21934 2144 21950 2208
rect 22014 2144 22030 2208
rect 22094 2144 22100 2208
rect 21784 2143 22100 2144
rect 28730 2208 29046 2209
rect 28730 2144 28736 2208
rect 28800 2144 28816 2208
rect 28880 2144 28896 2208
rect 28960 2144 28976 2208
rect 29040 2144 29046 2208
rect 28730 2143 29046 2144
rect 29200 2002 30000 2032
rect 24810 1942 30000 2002
rect 12750 1396 12756 1460
rect 12820 1458 12826 1460
rect 24810 1458 24870 1942
rect 29200 1912 30000 1942
rect 12820 1398 24870 1458
rect 12820 1396 12826 1398
<< via3 >>
rect 16436 31724 16500 31788
rect 7898 31580 7962 31584
rect 7898 31524 7902 31580
rect 7902 31524 7958 31580
rect 7958 31524 7962 31580
rect 7898 31520 7962 31524
rect 7978 31580 8042 31584
rect 7978 31524 7982 31580
rect 7982 31524 8038 31580
rect 8038 31524 8042 31580
rect 7978 31520 8042 31524
rect 8058 31580 8122 31584
rect 8058 31524 8062 31580
rect 8062 31524 8118 31580
rect 8118 31524 8122 31580
rect 8058 31520 8122 31524
rect 8138 31580 8202 31584
rect 8138 31524 8142 31580
rect 8142 31524 8198 31580
rect 8198 31524 8202 31580
rect 8138 31520 8202 31524
rect 14844 31580 14908 31584
rect 14844 31524 14848 31580
rect 14848 31524 14904 31580
rect 14904 31524 14908 31580
rect 14844 31520 14908 31524
rect 14924 31580 14988 31584
rect 14924 31524 14928 31580
rect 14928 31524 14984 31580
rect 14984 31524 14988 31580
rect 14924 31520 14988 31524
rect 15004 31580 15068 31584
rect 15004 31524 15008 31580
rect 15008 31524 15064 31580
rect 15064 31524 15068 31580
rect 15004 31520 15068 31524
rect 15084 31580 15148 31584
rect 15084 31524 15088 31580
rect 15088 31524 15144 31580
rect 15144 31524 15148 31580
rect 15084 31520 15148 31524
rect 21790 31580 21854 31584
rect 21790 31524 21794 31580
rect 21794 31524 21850 31580
rect 21850 31524 21854 31580
rect 21790 31520 21854 31524
rect 21870 31580 21934 31584
rect 21870 31524 21874 31580
rect 21874 31524 21930 31580
rect 21930 31524 21934 31580
rect 21870 31520 21934 31524
rect 21950 31580 22014 31584
rect 21950 31524 21954 31580
rect 21954 31524 22010 31580
rect 22010 31524 22014 31580
rect 21950 31520 22014 31524
rect 22030 31580 22094 31584
rect 22030 31524 22034 31580
rect 22034 31524 22090 31580
rect 22090 31524 22094 31580
rect 22030 31520 22094 31524
rect 28736 31580 28800 31584
rect 28736 31524 28740 31580
rect 28740 31524 28796 31580
rect 28796 31524 28800 31580
rect 28736 31520 28800 31524
rect 28816 31580 28880 31584
rect 28816 31524 28820 31580
rect 28820 31524 28876 31580
rect 28876 31524 28880 31580
rect 28816 31520 28880 31524
rect 28896 31580 28960 31584
rect 28896 31524 28900 31580
rect 28900 31524 28956 31580
rect 28956 31524 28960 31580
rect 28896 31520 28960 31524
rect 28976 31580 29040 31584
rect 28976 31524 28980 31580
rect 28980 31524 29036 31580
rect 29036 31524 29040 31580
rect 28976 31520 29040 31524
rect 15332 31316 15396 31380
rect 4425 31036 4489 31040
rect 4425 30980 4429 31036
rect 4429 30980 4485 31036
rect 4485 30980 4489 31036
rect 4425 30976 4489 30980
rect 4505 31036 4569 31040
rect 4505 30980 4509 31036
rect 4509 30980 4565 31036
rect 4565 30980 4569 31036
rect 4505 30976 4569 30980
rect 4585 31036 4649 31040
rect 4585 30980 4589 31036
rect 4589 30980 4645 31036
rect 4645 30980 4649 31036
rect 4585 30976 4649 30980
rect 4665 31036 4729 31040
rect 4665 30980 4669 31036
rect 4669 30980 4725 31036
rect 4725 30980 4729 31036
rect 4665 30976 4729 30980
rect 11371 31036 11435 31040
rect 11371 30980 11375 31036
rect 11375 30980 11431 31036
rect 11431 30980 11435 31036
rect 11371 30976 11435 30980
rect 11451 31036 11515 31040
rect 11451 30980 11455 31036
rect 11455 30980 11511 31036
rect 11511 30980 11515 31036
rect 11451 30976 11515 30980
rect 11531 31036 11595 31040
rect 11531 30980 11535 31036
rect 11535 30980 11591 31036
rect 11591 30980 11595 31036
rect 11531 30976 11595 30980
rect 11611 31036 11675 31040
rect 11611 30980 11615 31036
rect 11615 30980 11671 31036
rect 11671 30980 11675 31036
rect 11611 30976 11675 30980
rect 18317 31036 18381 31040
rect 18317 30980 18321 31036
rect 18321 30980 18377 31036
rect 18377 30980 18381 31036
rect 18317 30976 18381 30980
rect 18397 31036 18461 31040
rect 18397 30980 18401 31036
rect 18401 30980 18457 31036
rect 18457 30980 18461 31036
rect 18397 30976 18461 30980
rect 18477 31036 18541 31040
rect 18477 30980 18481 31036
rect 18481 30980 18537 31036
rect 18537 30980 18541 31036
rect 18477 30976 18541 30980
rect 18557 31036 18621 31040
rect 18557 30980 18561 31036
rect 18561 30980 18617 31036
rect 18617 30980 18621 31036
rect 18557 30976 18621 30980
rect 25263 31036 25327 31040
rect 25263 30980 25267 31036
rect 25267 30980 25323 31036
rect 25323 30980 25327 31036
rect 25263 30976 25327 30980
rect 25343 31036 25407 31040
rect 25343 30980 25347 31036
rect 25347 30980 25403 31036
rect 25403 30980 25407 31036
rect 25343 30976 25407 30980
rect 25423 31036 25487 31040
rect 25423 30980 25427 31036
rect 25427 30980 25483 31036
rect 25483 30980 25487 31036
rect 25423 30976 25487 30980
rect 25503 31036 25567 31040
rect 25503 30980 25507 31036
rect 25507 30980 25563 31036
rect 25563 30980 25567 31036
rect 25503 30976 25567 30980
rect 7898 30492 7962 30496
rect 7898 30436 7902 30492
rect 7902 30436 7958 30492
rect 7958 30436 7962 30492
rect 7898 30432 7962 30436
rect 7978 30492 8042 30496
rect 7978 30436 7982 30492
rect 7982 30436 8038 30492
rect 8038 30436 8042 30492
rect 7978 30432 8042 30436
rect 8058 30492 8122 30496
rect 8058 30436 8062 30492
rect 8062 30436 8118 30492
rect 8118 30436 8122 30492
rect 8058 30432 8122 30436
rect 8138 30492 8202 30496
rect 8138 30436 8142 30492
rect 8142 30436 8198 30492
rect 8198 30436 8202 30492
rect 8138 30432 8202 30436
rect 14844 30492 14908 30496
rect 14844 30436 14848 30492
rect 14848 30436 14904 30492
rect 14904 30436 14908 30492
rect 14844 30432 14908 30436
rect 14924 30492 14988 30496
rect 14924 30436 14928 30492
rect 14928 30436 14984 30492
rect 14984 30436 14988 30492
rect 14924 30432 14988 30436
rect 15004 30492 15068 30496
rect 15004 30436 15008 30492
rect 15008 30436 15064 30492
rect 15064 30436 15068 30492
rect 15004 30432 15068 30436
rect 15084 30492 15148 30496
rect 15084 30436 15088 30492
rect 15088 30436 15144 30492
rect 15144 30436 15148 30492
rect 15084 30432 15148 30436
rect 21790 30492 21854 30496
rect 21790 30436 21794 30492
rect 21794 30436 21850 30492
rect 21850 30436 21854 30492
rect 21790 30432 21854 30436
rect 21870 30492 21934 30496
rect 21870 30436 21874 30492
rect 21874 30436 21930 30492
rect 21930 30436 21934 30492
rect 21870 30432 21934 30436
rect 21950 30492 22014 30496
rect 21950 30436 21954 30492
rect 21954 30436 22010 30492
rect 22010 30436 22014 30492
rect 21950 30432 22014 30436
rect 22030 30492 22094 30496
rect 22030 30436 22034 30492
rect 22034 30436 22090 30492
rect 22090 30436 22094 30492
rect 22030 30432 22094 30436
rect 28736 30492 28800 30496
rect 28736 30436 28740 30492
rect 28740 30436 28796 30492
rect 28796 30436 28800 30492
rect 28736 30432 28800 30436
rect 28816 30492 28880 30496
rect 28816 30436 28820 30492
rect 28820 30436 28876 30492
rect 28876 30436 28880 30492
rect 28816 30432 28880 30436
rect 28896 30492 28960 30496
rect 28896 30436 28900 30492
rect 28900 30436 28956 30492
rect 28956 30436 28960 30492
rect 28896 30432 28960 30436
rect 28976 30492 29040 30496
rect 28976 30436 28980 30492
rect 28980 30436 29036 30492
rect 29036 30436 29040 30492
rect 28976 30432 29040 30436
rect 6868 30364 6932 30428
rect 16620 30364 16684 30428
rect 14596 30092 14660 30156
rect 4425 29948 4489 29952
rect 4425 29892 4429 29948
rect 4429 29892 4485 29948
rect 4485 29892 4489 29948
rect 4425 29888 4489 29892
rect 4505 29948 4569 29952
rect 4505 29892 4509 29948
rect 4509 29892 4565 29948
rect 4565 29892 4569 29948
rect 4505 29888 4569 29892
rect 4585 29948 4649 29952
rect 4585 29892 4589 29948
rect 4589 29892 4645 29948
rect 4645 29892 4649 29948
rect 4585 29888 4649 29892
rect 4665 29948 4729 29952
rect 4665 29892 4669 29948
rect 4669 29892 4725 29948
rect 4725 29892 4729 29948
rect 4665 29888 4729 29892
rect 11371 29948 11435 29952
rect 11371 29892 11375 29948
rect 11375 29892 11431 29948
rect 11431 29892 11435 29948
rect 11371 29888 11435 29892
rect 11451 29948 11515 29952
rect 11451 29892 11455 29948
rect 11455 29892 11511 29948
rect 11511 29892 11515 29948
rect 11451 29888 11515 29892
rect 11531 29948 11595 29952
rect 11531 29892 11535 29948
rect 11535 29892 11591 29948
rect 11591 29892 11595 29948
rect 11531 29888 11595 29892
rect 11611 29948 11675 29952
rect 11611 29892 11615 29948
rect 11615 29892 11671 29948
rect 11671 29892 11675 29948
rect 11611 29888 11675 29892
rect 18317 29948 18381 29952
rect 18317 29892 18321 29948
rect 18321 29892 18377 29948
rect 18377 29892 18381 29948
rect 18317 29888 18381 29892
rect 18397 29948 18461 29952
rect 18397 29892 18401 29948
rect 18401 29892 18457 29948
rect 18457 29892 18461 29948
rect 18397 29888 18461 29892
rect 18477 29948 18541 29952
rect 18477 29892 18481 29948
rect 18481 29892 18537 29948
rect 18537 29892 18541 29948
rect 18477 29888 18541 29892
rect 18557 29948 18621 29952
rect 18557 29892 18561 29948
rect 18561 29892 18617 29948
rect 18617 29892 18621 29948
rect 18557 29888 18621 29892
rect 25263 29948 25327 29952
rect 25263 29892 25267 29948
rect 25267 29892 25323 29948
rect 25323 29892 25327 29948
rect 25263 29888 25327 29892
rect 25343 29948 25407 29952
rect 25343 29892 25347 29948
rect 25347 29892 25403 29948
rect 25403 29892 25407 29948
rect 25343 29888 25407 29892
rect 25423 29948 25487 29952
rect 25423 29892 25427 29948
rect 25427 29892 25483 29948
rect 25483 29892 25487 29948
rect 25423 29888 25487 29892
rect 25503 29948 25567 29952
rect 25503 29892 25507 29948
rect 25507 29892 25563 29948
rect 25563 29892 25567 29948
rect 25503 29888 25567 29892
rect 15332 29684 15396 29748
rect 15700 29684 15764 29748
rect 12940 29548 13004 29612
rect 16620 29472 16684 29476
rect 16620 29416 16670 29472
rect 16670 29416 16684 29472
rect 16620 29412 16684 29416
rect 7898 29404 7962 29408
rect 7898 29348 7902 29404
rect 7902 29348 7958 29404
rect 7958 29348 7962 29404
rect 7898 29344 7962 29348
rect 7978 29404 8042 29408
rect 7978 29348 7982 29404
rect 7982 29348 8038 29404
rect 8038 29348 8042 29404
rect 7978 29344 8042 29348
rect 8058 29404 8122 29408
rect 8058 29348 8062 29404
rect 8062 29348 8118 29404
rect 8118 29348 8122 29404
rect 8058 29344 8122 29348
rect 8138 29404 8202 29408
rect 8138 29348 8142 29404
rect 8142 29348 8198 29404
rect 8198 29348 8202 29404
rect 8138 29344 8202 29348
rect 14844 29404 14908 29408
rect 14844 29348 14848 29404
rect 14848 29348 14904 29404
rect 14904 29348 14908 29404
rect 14844 29344 14908 29348
rect 14924 29404 14988 29408
rect 14924 29348 14928 29404
rect 14928 29348 14984 29404
rect 14984 29348 14988 29404
rect 14924 29344 14988 29348
rect 15004 29404 15068 29408
rect 15004 29348 15008 29404
rect 15008 29348 15064 29404
rect 15064 29348 15068 29404
rect 15004 29344 15068 29348
rect 15084 29404 15148 29408
rect 15084 29348 15088 29404
rect 15088 29348 15144 29404
rect 15144 29348 15148 29404
rect 15084 29344 15148 29348
rect 21790 29404 21854 29408
rect 21790 29348 21794 29404
rect 21794 29348 21850 29404
rect 21850 29348 21854 29404
rect 21790 29344 21854 29348
rect 21870 29404 21934 29408
rect 21870 29348 21874 29404
rect 21874 29348 21930 29404
rect 21930 29348 21934 29404
rect 21870 29344 21934 29348
rect 21950 29404 22014 29408
rect 21950 29348 21954 29404
rect 21954 29348 22010 29404
rect 22010 29348 22014 29404
rect 21950 29344 22014 29348
rect 22030 29404 22094 29408
rect 22030 29348 22034 29404
rect 22034 29348 22090 29404
rect 22090 29348 22094 29404
rect 22030 29344 22094 29348
rect 28736 29404 28800 29408
rect 28736 29348 28740 29404
rect 28740 29348 28796 29404
rect 28796 29348 28800 29404
rect 28736 29344 28800 29348
rect 28816 29404 28880 29408
rect 28816 29348 28820 29404
rect 28820 29348 28876 29404
rect 28876 29348 28880 29404
rect 28816 29344 28880 29348
rect 28896 29404 28960 29408
rect 28896 29348 28900 29404
rect 28900 29348 28956 29404
rect 28956 29348 28960 29404
rect 28896 29344 28960 29348
rect 28976 29404 29040 29408
rect 28976 29348 28980 29404
rect 28980 29348 29036 29404
rect 29036 29348 29040 29404
rect 28976 29344 29040 29348
rect 15700 29140 15764 29204
rect 16436 29140 16500 29204
rect 4425 28860 4489 28864
rect 4425 28804 4429 28860
rect 4429 28804 4485 28860
rect 4485 28804 4489 28860
rect 4425 28800 4489 28804
rect 4505 28860 4569 28864
rect 4505 28804 4509 28860
rect 4509 28804 4565 28860
rect 4565 28804 4569 28860
rect 4505 28800 4569 28804
rect 4585 28860 4649 28864
rect 4585 28804 4589 28860
rect 4589 28804 4645 28860
rect 4645 28804 4649 28860
rect 4585 28800 4649 28804
rect 4665 28860 4729 28864
rect 4665 28804 4669 28860
rect 4669 28804 4725 28860
rect 4725 28804 4729 28860
rect 4665 28800 4729 28804
rect 11371 28860 11435 28864
rect 11371 28804 11375 28860
rect 11375 28804 11431 28860
rect 11431 28804 11435 28860
rect 11371 28800 11435 28804
rect 11451 28860 11515 28864
rect 11451 28804 11455 28860
rect 11455 28804 11511 28860
rect 11511 28804 11515 28860
rect 11451 28800 11515 28804
rect 11531 28860 11595 28864
rect 11531 28804 11535 28860
rect 11535 28804 11591 28860
rect 11591 28804 11595 28860
rect 11531 28800 11595 28804
rect 11611 28860 11675 28864
rect 11611 28804 11615 28860
rect 11615 28804 11671 28860
rect 11671 28804 11675 28860
rect 11611 28800 11675 28804
rect 18317 28860 18381 28864
rect 18317 28804 18321 28860
rect 18321 28804 18377 28860
rect 18377 28804 18381 28860
rect 18317 28800 18381 28804
rect 18397 28860 18461 28864
rect 18397 28804 18401 28860
rect 18401 28804 18457 28860
rect 18457 28804 18461 28860
rect 18397 28800 18461 28804
rect 18477 28860 18541 28864
rect 18477 28804 18481 28860
rect 18481 28804 18537 28860
rect 18537 28804 18541 28860
rect 18477 28800 18541 28804
rect 18557 28860 18621 28864
rect 18557 28804 18561 28860
rect 18561 28804 18617 28860
rect 18617 28804 18621 28860
rect 18557 28800 18621 28804
rect 25263 28860 25327 28864
rect 25263 28804 25267 28860
rect 25267 28804 25323 28860
rect 25323 28804 25327 28860
rect 25263 28800 25327 28804
rect 25343 28860 25407 28864
rect 25343 28804 25347 28860
rect 25347 28804 25403 28860
rect 25403 28804 25407 28860
rect 25343 28800 25407 28804
rect 25423 28860 25487 28864
rect 25423 28804 25427 28860
rect 25427 28804 25483 28860
rect 25483 28804 25487 28860
rect 25423 28800 25487 28804
rect 25503 28860 25567 28864
rect 25503 28804 25507 28860
rect 25507 28804 25563 28860
rect 25563 28804 25567 28860
rect 25503 28800 25567 28804
rect 7898 28316 7962 28320
rect 7898 28260 7902 28316
rect 7902 28260 7958 28316
rect 7958 28260 7962 28316
rect 7898 28256 7962 28260
rect 7978 28316 8042 28320
rect 7978 28260 7982 28316
rect 7982 28260 8038 28316
rect 8038 28260 8042 28316
rect 7978 28256 8042 28260
rect 8058 28316 8122 28320
rect 8058 28260 8062 28316
rect 8062 28260 8118 28316
rect 8118 28260 8122 28316
rect 8058 28256 8122 28260
rect 8138 28316 8202 28320
rect 8138 28260 8142 28316
rect 8142 28260 8198 28316
rect 8198 28260 8202 28316
rect 8138 28256 8202 28260
rect 14844 28316 14908 28320
rect 14844 28260 14848 28316
rect 14848 28260 14904 28316
rect 14904 28260 14908 28316
rect 14844 28256 14908 28260
rect 14924 28316 14988 28320
rect 14924 28260 14928 28316
rect 14928 28260 14984 28316
rect 14984 28260 14988 28316
rect 14924 28256 14988 28260
rect 15004 28316 15068 28320
rect 15004 28260 15008 28316
rect 15008 28260 15064 28316
rect 15064 28260 15068 28316
rect 15004 28256 15068 28260
rect 15084 28316 15148 28320
rect 15084 28260 15088 28316
rect 15088 28260 15144 28316
rect 15144 28260 15148 28316
rect 15084 28256 15148 28260
rect 21790 28316 21854 28320
rect 21790 28260 21794 28316
rect 21794 28260 21850 28316
rect 21850 28260 21854 28316
rect 21790 28256 21854 28260
rect 21870 28316 21934 28320
rect 21870 28260 21874 28316
rect 21874 28260 21930 28316
rect 21930 28260 21934 28316
rect 21870 28256 21934 28260
rect 21950 28316 22014 28320
rect 21950 28260 21954 28316
rect 21954 28260 22010 28316
rect 22010 28260 22014 28316
rect 21950 28256 22014 28260
rect 22030 28316 22094 28320
rect 22030 28260 22034 28316
rect 22034 28260 22090 28316
rect 22090 28260 22094 28316
rect 22030 28256 22094 28260
rect 28736 28316 28800 28320
rect 28736 28260 28740 28316
rect 28740 28260 28796 28316
rect 28796 28260 28800 28316
rect 28736 28256 28800 28260
rect 28816 28316 28880 28320
rect 28816 28260 28820 28316
rect 28820 28260 28876 28316
rect 28876 28260 28880 28316
rect 28816 28256 28880 28260
rect 28896 28316 28960 28320
rect 28896 28260 28900 28316
rect 28900 28260 28956 28316
rect 28956 28260 28960 28316
rect 28896 28256 28960 28260
rect 28976 28316 29040 28320
rect 28976 28260 28980 28316
rect 28980 28260 29036 28316
rect 29036 28260 29040 28316
rect 28976 28256 29040 28260
rect 4425 27772 4489 27776
rect 4425 27716 4429 27772
rect 4429 27716 4485 27772
rect 4485 27716 4489 27772
rect 4425 27712 4489 27716
rect 4505 27772 4569 27776
rect 4505 27716 4509 27772
rect 4509 27716 4565 27772
rect 4565 27716 4569 27772
rect 4505 27712 4569 27716
rect 4585 27772 4649 27776
rect 4585 27716 4589 27772
rect 4589 27716 4645 27772
rect 4645 27716 4649 27772
rect 4585 27712 4649 27716
rect 4665 27772 4729 27776
rect 4665 27716 4669 27772
rect 4669 27716 4725 27772
rect 4725 27716 4729 27772
rect 4665 27712 4729 27716
rect 11371 27772 11435 27776
rect 11371 27716 11375 27772
rect 11375 27716 11431 27772
rect 11431 27716 11435 27772
rect 11371 27712 11435 27716
rect 11451 27772 11515 27776
rect 11451 27716 11455 27772
rect 11455 27716 11511 27772
rect 11511 27716 11515 27772
rect 11451 27712 11515 27716
rect 11531 27772 11595 27776
rect 11531 27716 11535 27772
rect 11535 27716 11591 27772
rect 11591 27716 11595 27772
rect 11531 27712 11595 27716
rect 11611 27772 11675 27776
rect 11611 27716 11615 27772
rect 11615 27716 11671 27772
rect 11671 27716 11675 27772
rect 11611 27712 11675 27716
rect 12756 27916 12820 27980
rect 18317 27772 18381 27776
rect 18317 27716 18321 27772
rect 18321 27716 18377 27772
rect 18377 27716 18381 27772
rect 18317 27712 18381 27716
rect 18397 27772 18461 27776
rect 18397 27716 18401 27772
rect 18401 27716 18457 27772
rect 18457 27716 18461 27772
rect 18397 27712 18461 27716
rect 18477 27772 18541 27776
rect 18477 27716 18481 27772
rect 18481 27716 18537 27772
rect 18537 27716 18541 27772
rect 18477 27712 18541 27716
rect 18557 27772 18621 27776
rect 18557 27716 18561 27772
rect 18561 27716 18617 27772
rect 18617 27716 18621 27772
rect 18557 27712 18621 27716
rect 25263 27772 25327 27776
rect 25263 27716 25267 27772
rect 25267 27716 25323 27772
rect 25323 27716 25327 27772
rect 25263 27712 25327 27716
rect 25343 27772 25407 27776
rect 25343 27716 25347 27772
rect 25347 27716 25403 27772
rect 25403 27716 25407 27772
rect 25343 27712 25407 27716
rect 25423 27772 25487 27776
rect 25423 27716 25427 27772
rect 25427 27716 25483 27772
rect 25483 27716 25487 27772
rect 25423 27712 25487 27716
rect 25503 27772 25567 27776
rect 25503 27716 25507 27772
rect 25507 27716 25563 27772
rect 25563 27716 25567 27772
rect 25503 27712 25567 27716
rect 6868 27372 6932 27436
rect 7898 27228 7962 27232
rect 7898 27172 7902 27228
rect 7902 27172 7958 27228
rect 7958 27172 7962 27228
rect 7898 27168 7962 27172
rect 7978 27228 8042 27232
rect 7978 27172 7982 27228
rect 7982 27172 8038 27228
rect 8038 27172 8042 27228
rect 7978 27168 8042 27172
rect 8058 27228 8122 27232
rect 8058 27172 8062 27228
rect 8062 27172 8118 27228
rect 8118 27172 8122 27228
rect 8058 27168 8122 27172
rect 8138 27228 8202 27232
rect 8138 27172 8142 27228
rect 8142 27172 8198 27228
rect 8198 27172 8202 27228
rect 8138 27168 8202 27172
rect 12940 27296 13004 27300
rect 12940 27240 12990 27296
rect 12990 27240 13004 27296
rect 12940 27236 13004 27240
rect 14844 27228 14908 27232
rect 14844 27172 14848 27228
rect 14848 27172 14904 27228
rect 14904 27172 14908 27228
rect 14844 27168 14908 27172
rect 14924 27228 14988 27232
rect 14924 27172 14928 27228
rect 14928 27172 14984 27228
rect 14984 27172 14988 27228
rect 14924 27168 14988 27172
rect 15004 27228 15068 27232
rect 15004 27172 15008 27228
rect 15008 27172 15064 27228
rect 15064 27172 15068 27228
rect 15004 27168 15068 27172
rect 15084 27228 15148 27232
rect 15084 27172 15088 27228
rect 15088 27172 15144 27228
rect 15144 27172 15148 27228
rect 15084 27168 15148 27172
rect 21790 27228 21854 27232
rect 21790 27172 21794 27228
rect 21794 27172 21850 27228
rect 21850 27172 21854 27228
rect 21790 27168 21854 27172
rect 21870 27228 21934 27232
rect 21870 27172 21874 27228
rect 21874 27172 21930 27228
rect 21930 27172 21934 27228
rect 21870 27168 21934 27172
rect 21950 27228 22014 27232
rect 21950 27172 21954 27228
rect 21954 27172 22010 27228
rect 22010 27172 22014 27228
rect 21950 27168 22014 27172
rect 22030 27228 22094 27232
rect 22030 27172 22034 27228
rect 22034 27172 22090 27228
rect 22090 27172 22094 27228
rect 22030 27168 22094 27172
rect 28736 27228 28800 27232
rect 28736 27172 28740 27228
rect 28740 27172 28796 27228
rect 28796 27172 28800 27228
rect 28736 27168 28800 27172
rect 28816 27228 28880 27232
rect 28816 27172 28820 27228
rect 28820 27172 28876 27228
rect 28876 27172 28880 27228
rect 28816 27168 28880 27172
rect 28896 27228 28960 27232
rect 28896 27172 28900 27228
rect 28900 27172 28956 27228
rect 28956 27172 28960 27228
rect 28896 27168 28960 27172
rect 28976 27228 29040 27232
rect 28976 27172 28980 27228
rect 28980 27172 29036 27228
rect 29036 27172 29040 27228
rect 28976 27168 29040 27172
rect 4425 26684 4489 26688
rect 4425 26628 4429 26684
rect 4429 26628 4485 26684
rect 4485 26628 4489 26684
rect 4425 26624 4489 26628
rect 4505 26684 4569 26688
rect 4505 26628 4509 26684
rect 4509 26628 4565 26684
rect 4565 26628 4569 26684
rect 4505 26624 4569 26628
rect 4585 26684 4649 26688
rect 4585 26628 4589 26684
rect 4589 26628 4645 26684
rect 4645 26628 4649 26684
rect 4585 26624 4649 26628
rect 4665 26684 4729 26688
rect 4665 26628 4669 26684
rect 4669 26628 4725 26684
rect 4725 26628 4729 26684
rect 4665 26624 4729 26628
rect 11371 26684 11435 26688
rect 11371 26628 11375 26684
rect 11375 26628 11431 26684
rect 11431 26628 11435 26684
rect 11371 26624 11435 26628
rect 11451 26684 11515 26688
rect 11451 26628 11455 26684
rect 11455 26628 11511 26684
rect 11511 26628 11515 26684
rect 11451 26624 11515 26628
rect 11531 26684 11595 26688
rect 11531 26628 11535 26684
rect 11535 26628 11591 26684
rect 11591 26628 11595 26684
rect 11531 26624 11595 26628
rect 11611 26684 11675 26688
rect 11611 26628 11615 26684
rect 11615 26628 11671 26684
rect 11671 26628 11675 26684
rect 11611 26624 11675 26628
rect 18317 26684 18381 26688
rect 18317 26628 18321 26684
rect 18321 26628 18377 26684
rect 18377 26628 18381 26684
rect 18317 26624 18381 26628
rect 18397 26684 18461 26688
rect 18397 26628 18401 26684
rect 18401 26628 18457 26684
rect 18457 26628 18461 26684
rect 18397 26624 18461 26628
rect 18477 26684 18541 26688
rect 18477 26628 18481 26684
rect 18481 26628 18537 26684
rect 18537 26628 18541 26684
rect 18477 26624 18541 26628
rect 18557 26684 18621 26688
rect 18557 26628 18561 26684
rect 18561 26628 18617 26684
rect 18617 26628 18621 26684
rect 18557 26624 18621 26628
rect 25263 26684 25327 26688
rect 25263 26628 25267 26684
rect 25267 26628 25323 26684
rect 25323 26628 25327 26684
rect 25263 26624 25327 26628
rect 25343 26684 25407 26688
rect 25343 26628 25347 26684
rect 25347 26628 25403 26684
rect 25403 26628 25407 26684
rect 25343 26624 25407 26628
rect 25423 26684 25487 26688
rect 25423 26628 25427 26684
rect 25427 26628 25483 26684
rect 25483 26628 25487 26684
rect 25423 26624 25487 26628
rect 25503 26684 25567 26688
rect 25503 26628 25507 26684
rect 25507 26628 25563 26684
rect 25563 26628 25567 26684
rect 25503 26624 25567 26628
rect 14596 26420 14660 26484
rect 7898 26140 7962 26144
rect 7898 26084 7902 26140
rect 7902 26084 7958 26140
rect 7958 26084 7962 26140
rect 7898 26080 7962 26084
rect 7978 26140 8042 26144
rect 7978 26084 7982 26140
rect 7982 26084 8038 26140
rect 8038 26084 8042 26140
rect 7978 26080 8042 26084
rect 8058 26140 8122 26144
rect 8058 26084 8062 26140
rect 8062 26084 8118 26140
rect 8118 26084 8122 26140
rect 8058 26080 8122 26084
rect 8138 26140 8202 26144
rect 8138 26084 8142 26140
rect 8142 26084 8198 26140
rect 8198 26084 8202 26140
rect 8138 26080 8202 26084
rect 14844 26140 14908 26144
rect 14844 26084 14848 26140
rect 14848 26084 14904 26140
rect 14904 26084 14908 26140
rect 14844 26080 14908 26084
rect 14924 26140 14988 26144
rect 14924 26084 14928 26140
rect 14928 26084 14984 26140
rect 14984 26084 14988 26140
rect 14924 26080 14988 26084
rect 15004 26140 15068 26144
rect 15004 26084 15008 26140
rect 15008 26084 15064 26140
rect 15064 26084 15068 26140
rect 15004 26080 15068 26084
rect 15084 26140 15148 26144
rect 15084 26084 15088 26140
rect 15088 26084 15144 26140
rect 15144 26084 15148 26140
rect 15084 26080 15148 26084
rect 21790 26140 21854 26144
rect 21790 26084 21794 26140
rect 21794 26084 21850 26140
rect 21850 26084 21854 26140
rect 21790 26080 21854 26084
rect 21870 26140 21934 26144
rect 21870 26084 21874 26140
rect 21874 26084 21930 26140
rect 21930 26084 21934 26140
rect 21870 26080 21934 26084
rect 21950 26140 22014 26144
rect 21950 26084 21954 26140
rect 21954 26084 22010 26140
rect 22010 26084 22014 26140
rect 21950 26080 22014 26084
rect 22030 26140 22094 26144
rect 22030 26084 22034 26140
rect 22034 26084 22090 26140
rect 22090 26084 22094 26140
rect 22030 26080 22094 26084
rect 28736 26140 28800 26144
rect 28736 26084 28740 26140
rect 28740 26084 28796 26140
rect 28796 26084 28800 26140
rect 28736 26080 28800 26084
rect 28816 26140 28880 26144
rect 28816 26084 28820 26140
rect 28820 26084 28876 26140
rect 28876 26084 28880 26140
rect 28816 26080 28880 26084
rect 28896 26140 28960 26144
rect 28896 26084 28900 26140
rect 28900 26084 28956 26140
rect 28956 26084 28960 26140
rect 28896 26080 28960 26084
rect 28976 26140 29040 26144
rect 28976 26084 28980 26140
rect 28980 26084 29036 26140
rect 29036 26084 29040 26140
rect 28976 26080 29040 26084
rect 4425 25596 4489 25600
rect 4425 25540 4429 25596
rect 4429 25540 4485 25596
rect 4485 25540 4489 25596
rect 4425 25536 4489 25540
rect 4505 25596 4569 25600
rect 4505 25540 4509 25596
rect 4509 25540 4565 25596
rect 4565 25540 4569 25596
rect 4505 25536 4569 25540
rect 4585 25596 4649 25600
rect 4585 25540 4589 25596
rect 4589 25540 4645 25596
rect 4645 25540 4649 25596
rect 4585 25536 4649 25540
rect 4665 25596 4729 25600
rect 4665 25540 4669 25596
rect 4669 25540 4725 25596
rect 4725 25540 4729 25596
rect 4665 25536 4729 25540
rect 11371 25596 11435 25600
rect 11371 25540 11375 25596
rect 11375 25540 11431 25596
rect 11431 25540 11435 25596
rect 11371 25536 11435 25540
rect 11451 25596 11515 25600
rect 11451 25540 11455 25596
rect 11455 25540 11511 25596
rect 11511 25540 11515 25596
rect 11451 25536 11515 25540
rect 11531 25596 11595 25600
rect 11531 25540 11535 25596
rect 11535 25540 11591 25596
rect 11591 25540 11595 25596
rect 11531 25536 11595 25540
rect 11611 25596 11675 25600
rect 11611 25540 11615 25596
rect 11615 25540 11671 25596
rect 11671 25540 11675 25596
rect 11611 25536 11675 25540
rect 18317 25596 18381 25600
rect 18317 25540 18321 25596
rect 18321 25540 18377 25596
rect 18377 25540 18381 25596
rect 18317 25536 18381 25540
rect 18397 25596 18461 25600
rect 18397 25540 18401 25596
rect 18401 25540 18457 25596
rect 18457 25540 18461 25596
rect 18397 25536 18461 25540
rect 18477 25596 18541 25600
rect 18477 25540 18481 25596
rect 18481 25540 18537 25596
rect 18537 25540 18541 25596
rect 18477 25536 18541 25540
rect 18557 25596 18621 25600
rect 18557 25540 18561 25596
rect 18561 25540 18617 25596
rect 18617 25540 18621 25596
rect 18557 25536 18621 25540
rect 25263 25596 25327 25600
rect 25263 25540 25267 25596
rect 25267 25540 25323 25596
rect 25323 25540 25327 25596
rect 25263 25536 25327 25540
rect 25343 25596 25407 25600
rect 25343 25540 25347 25596
rect 25347 25540 25403 25596
rect 25403 25540 25407 25596
rect 25343 25536 25407 25540
rect 25423 25596 25487 25600
rect 25423 25540 25427 25596
rect 25427 25540 25483 25596
rect 25483 25540 25487 25596
rect 25423 25536 25487 25540
rect 25503 25596 25567 25600
rect 25503 25540 25507 25596
rect 25507 25540 25563 25596
rect 25563 25540 25567 25596
rect 25503 25536 25567 25540
rect 7898 25052 7962 25056
rect 7898 24996 7902 25052
rect 7902 24996 7958 25052
rect 7958 24996 7962 25052
rect 7898 24992 7962 24996
rect 7978 25052 8042 25056
rect 7978 24996 7982 25052
rect 7982 24996 8038 25052
rect 8038 24996 8042 25052
rect 7978 24992 8042 24996
rect 8058 25052 8122 25056
rect 8058 24996 8062 25052
rect 8062 24996 8118 25052
rect 8118 24996 8122 25052
rect 8058 24992 8122 24996
rect 8138 25052 8202 25056
rect 8138 24996 8142 25052
rect 8142 24996 8198 25052
rect 8198 24996 8202 25052
rect 8138 24992 8202 24996
rect 14844 25052 14908 25056
rect 14844 24996 14848 25052
rect 14848 24996 14904 25052
rect 14904 24996 14908 25052
rect 14844 24992 14908 24996
rect 14924 25052 14988 25056
rect 14924 24996 14928 25052
rect 14928 24996 14984 25052
rect 14984 24996 14988 25052
rect 14924 24992 14988 24996
rect 15004 25052 15068 25056
rect 15004 24996 15008 25052
rect 15008 24996 15064 25052
rect 15064 24996 15068 25052
rect 15004 24992 15068 24996
rect 15084 25052 15148 25056
rect 15084 24996 15088 25052
rect 15088 24996 15144 25052
rect 15144 24996 15148 25052
rect 15084 24992 15148 24996
rect 21790 25052 21854 25056
rect 21790 24996 21794 25052
rect 21794 24996 21850 25052
rect 21850 24996 21854 25052
rect 21790 24992 21854 24996
rect 21870 25052 21934 25056
rect 21870 24996 21874 25052
rect 21874 24996 21930 25052
rect 21930 24996 21934 25052
rect 21870 24992 21934 24996
rect 21950 25052 22014 25056
rect 21950 24996 21954 25052
rect 21954 24996 22010 25052
rect 22010 24996 22014 25052
rect 21950 24992 22014 24996
rect 22030 25052 22094 25056
rect 22030 24996 22034 25052
rect 22034 24996 22090 25052
rect 22090 24996 22094 25052
rect 22030 24992 22094 24996
rect 28736 25052 28800 25056
rect 28736 24996 28740 25052
rect 28740 24996 28796 25052
rect 28796 24996 28800 25052
rect 28736 24992 28800 24996
rect 28816 25052 28880 25056
rect 28816 24996 28820 25052
rect 28820 24996 28876 25052
rect 28876 24996 28880 25052
rect 28816 24992 28880 24996
rect 28896 25052 28960 25056
rect 28896 24996 28900 25052
rect 28900 24996 28956 25052
rect 28956 24996 28960 25052
rect 28896 24992 28960 24996
rect 28976 25052 29040 25056
rect 28976 24996 28980 25052
rect 28980 24996 29036 25052
rect 29036 24996 29040 25052
rect 28976 24992 29040 24996
rect 4425 24508 4489 24512
rect 4425 24452 4429 24508
rect 4429 24452 4485 24508
rect 4485 24452 4489 24508
rect 4425 24448 4489 24452
rect 4505 24508 4569 24512
rect 4505 24452 4509 24508
rect 4509 24452 4565 24508
rect 4565 24452 4569 24508
rect 4505 24448 4569 24452
rect 4585 24508 4649 24512
rect 4585 24452 4589 24508
rect 4589 24452 4645 24508
rect 4645 24452 4649 24508
rect 4585 24448 4649 24452
rect 4665 24508 4729 24512
rect 4665 24452 4669 24508
rect 4669 24452 4725 24508
rect 4725 24452 4729 24508
rect 4665 24448 4729 24452
rect 11371 24508 11435 24512
rect 11371 24452 11375 24508
rect 11375 24452 11431 24508
rect 11431 24452 11435 24508
rect 11371 24448 11435 24452
rect 11451 24508 11515 24512
rect 11451 24452 11455 24508
rect 11455 24452 11511 24508
rect 11511 24452 11515 24508
rect 11451 24448 11515 24452
rect 11531 24508 11595 24512
rect 11531 24452 11535 24508
rect 11535 24452 11591 24508
rect 11591 24452 11595 24508
rect 11531 24448 11595 24452
rect 11611 24508 11675 24512
rect 11611 24452 11615 24508
rect 11615 24452 11671 24508
rect 11671 24452 11675 24508
rect 11611 24448 11675 24452
rect 18317 24508 18381 24512
rect 18317 24452 18321 24508
rect 18321 24452 18377 24508
rect 18377 24452 18381 24508
rect 18317 24448 18381 24452
rect 18397 24508 18461 24512
rect 18397 24452 18401 24508
rect 18401 24452 18457 24508
rect 18457 24452 18461 24508
rect 18397 24448 18461 24452
rect 18477 24508 18541 24512
rect 18477 24452 18481 24508
rect 18481 24452 18537 24508
rect 18537 24452 18541 24508
rect 18477 24448 18541 24452
rect 18557 24508 18621 24512
rect 18557 24452 18561 24508
rect 18561 24452 18617 24508
rect 18617 24452 18621 24508
rect 18557 24448 18621 24452
rect 25263 24508 25327 24512
rect 25263 24452 25267 24508
rect 25267 24452 25323 24508
rect 25323 24452 25327 24508
rect 25263 24448 25327 24452
rect 25343 24508 25407 24512
rect 25343 24452 25347 24508
rect 25347 24452 25403 24508
rect 25403 24452 25407 24508
rect 25343 24448 25407 24452
rect 25423 24508 25487 24512
rect 25423 24452 25427 24508
rect 25427 24452 25483 24508
rect 25483 24452 25487 24508
rect 25423 24448 25487 24452
rect 25503 24508 25567 24512
rect 25503 24452 25507 24508
rect 25507 24452 25563 24508
rect 25563 24452 25567 24508
rect 25503 24448 25567 24452
rect 7898 23964 7962 23968
rect 7898 23908 7902 23964
rect 7902 23908 7958 23964
rect 7958 23908 7962 23964
rect 7898 23904 7962 23908
rect 7978 23964 8042 23968
rect 7978 23908 7982 23964
rect 7982 23908 8038 23964
rect 8038 23908 8042 23964
rect 7978 23904 8042 23908
rect 8058 23964 8122 23968
rect 8058 23908 8062 23964
rect 8062 23908 8118 23964
rect 8118 23908 8122 23964
rect 8058 23904 8122 23908
rect 8138 23964 8202 23968
rect 8138 23908 8142 23964
rect 8142 23908 8198 23964
rect 8198 23908 8202 23964
rect 8138 23904 8202 23908
rect 14844 23964 14908 23968
rect 14844 23908 14848 23964
rect 14848 23908 14904 23964
rect 14904 23908 14908 23964
rect 14844 23904 14908 23908
rect 14924 23964 14988 23968
rect 14924 23908 14928 23964
rect 14928 23908 14984 23964
rect 14984 23908 14988 23964
rect 14924 23904 14988 23908
rect 15004 23964 15068 23968
rect 15004 23908 15008 23964
rect 15008 23908 15064 23964
rect 15064 23908 15068 23964
rect 15004 23904 15068 23908
rect 15084 23964 15148 23968
rect 15084 23908 15088 23964
rect 15088 23908 15144 23964
rect 15144 23908 15148 23964
rect 15084 23904 15148 23908
rect 21790 23964 21854 23968
rect 21790 23908 21794 23964
rect 21794 23908 21850 23964
rect 21850 23908 21854 23964
rect 21790 23904 21854 23908
rect 21870 23964 21934 23968
rect 21870 23908 21874 23964
rect 21874 23908 21930 23964
rect 21930 23908 21934 23964
rect 21870 23904 21934 23908
rect 21950 23964 22014 23968
rect 21950 23908 21954 23964
rect 21954 23908 22010 23964
rect 22010 23908 22014 23964
rect 21950 23904 22014 23908
rect 22030 23964 22094 23968
rect 22030 23908 22034 23964
rect 22034 23908 22090 23964
rect 22090 23908 22094 23964
rect 22030 23904 22094 23908
rect 28736 23964 28800 23968
rect 28736 23908 28740 23964
rect 28740 23908 28796 23964
rect 28796 23908 28800 23964
rect 28736 23904 28800 23908
rect 28816 23964 28880 23968
rect 28816 23908 28820 23964
rect 28820 23908 28876 23964
rect 28876 23908 28880 23964
rect 28816 23904 28880 23908
rect 28896 23964 28960 23968
rect 28896 23908 28900 23964
rect 28900 23908 28956 23964
rect 28956 23908 28960 23964
rect 28896 23904 28960 23908
rect 28976 23964 29040 23968
rect 28976 23908 28980 23964
rect 28980 23908 29036 23964
rect 29036 23908 29040 23964
rect 28976 23904 29040 23908
rect 4425 23420 4489 23424
rect 4425 23364 4429 23420
rect 4429 23364 4485 23420
rect 4485 23364 4489 23420
rect 4425 23360 4489 23364
rect 4505 23420 4569 23424
rect 4505 23364 4509 23420
rect 4509 23364 4565 23420
rect 4565 23364 4569 23420
rect 4505 23360 4569 23364
rect 4585 23420 4649 23424
rect 4585 23364 4589 23420
rect 4589 23364 4645 23420
rect 4645 23364 4649 23420
rect 4585 23360 4649 23364
rect 4665 23420 4729 23424
rect 4665 23364 4669 23420
rect 4669 23364 4725 23420
rect 4725 23364 4729 23420
rect 4665 23360 4729 23364
rect 11371 23420 11435 23424
rect 11371 23364 11375 23420
rect 11375 23364 11431 23420
rect 11431 23364 11435 23420
rect 11371 23360 11435 23364
rect 11451 23420 11515 23424
rect 11451 23364 11455 23420
rect 11455 23364 11511 23420
rect 11511 23364 11515 23420
rect 11451 23360 11515 23364
rect 11531 23420 11595 23424
rect 11531 23364 11535 23420
rect 11535 23364 11591 23420
rect 11591 23364 11595 23420
rect 11531 23360 11595 23364
rect 11611 23420 11675 23424
rect 11611 23364 11615 23420
rect 11615 23364 11671 23420
rect 11671 23364 11675 23420
rect 11611 23360 11675 23364
rect 18317 23420 18381 23424
rect 18317 23364 18321 23420
rect 18321 23364 18377 23420
rect 18377 23364 18381 23420
rect 18317 23360 18381 23364
rect 18397 23420 18461 23424
rect 18397 23364 18401 23420
rect 18401 23364 18457 23420
rect 18457 23364 18461 23420
rect 18397 23360 18461 23364
rect 18477 23420 18541 23424
rect 18477 23364 18481 23420
rect 18481 23364 18537 23420
rect 18537 23364 18541 23420
rect 18477 23360 18541 23364
rect 18557 23420 18621 23424
rect 18557 23364 18561 23420
rect 18561 23364 18617 23420
rect 18617 23364 18621 23420
rect 18557 23360 18621 23364
rect 25263 23420 25327 23424
rect 25263 23364 25267 23420
rect 25267 23364 25323 23420
rect 25323 23364 25327 23420
rect 25263 23360 25327 23364
rect 25343 23420 25407 23424
rect 25343 23364 25347 23420
rect 25347 23364 25403 23420
rect 25403 23364 25407 23420
rect 25343 23360 25407 23364
rect 25423 23420 25487 23424
rect 25423 23364 25427 23420
rect 25427 23364 25483 23420
rect 25483 23364 25487 23420
rect 25423 23360 25487 23364
rect 25503 23420 25567 23424
rect 25503 23364 25507 23420
rect 25507 23364 25563 23420
rect 25563 23364 25567 23420
rect 25503 23360 25567 23364
rect 7898 22876 7962 22880
rect 7898 22820 7902 22876
rect 7902 22820 7958 22876
rect 7958 22820 7962 22876
rect 7898 22816 7962 22820
rect 7978 22876 8042 22880
rect 7978 22820 7982 22876
rect 7982 22820 8038 22876
rect 8038 22820 8042 22876
rect 7978 22816 8042 22820
rect 8058 22876 8122 22880
rect 8058 22820 8062 22876
rect 8062 22820 8118 22876
rect 8118 22820 8122 22876
rect 8058 22816 8122 22820
rect 8138 22876 8202 22880
rect 8138 22820 8142 22876
rect 8142 22820 8198 22876
rect 8198 22820 8202 22876
rect 8138 22816 8202 22820
rect 14844 22876 14908 22880
rect 14844 22820 14848 22876
rect 14848 22820 14904 22876
rect 14904 22820 14908 22876
rect 14844 22816 14908 22820
rect 14924 22876 14988 22880
rect 14924 22820 14928 22876
rect 14928 22820 14984 22876
rect 14984 22820 14988 22876
rect 14924 22816 14988 22820
rect 15004 22876 15068 22880
rect 15004 22820 15008 22876
rect 15008 22820 15064 22876
rect 15064 22820 15068 22876
rect 15004 22816 15068 22820
rect 15084 22876 15148 22880
rect 15084 22820 15088 22876
rect 15088 22820 15144 22876
rect 15144 22820 15148 22876
rect 15084 22816 15148 22820
rect 21790 22876 21854 22880
rect 21790 22820 21794 22876
rect 21794 22820 21850 22876
rect 21850 22820 21854 22876
rect 21790 22816 21854 22820
rect 21870 22876 21934 22880
rect 21870 22820 21874 22876
rect 21874 22820 21930 22876
rect 21930 22820 21934 22876
rect 21870 22816 21934 22820
rect 21950 22876 22014 22880
rect 21950 22820 21954 22876
rect 21954 22820 22010 22876
rect 22010 22820 22014 22876
rect 21950 22816 22014 22820
rect 22030 22876 22094 22880
rect 22030 22820 22034 22876
rect 22034 22820 22090 22876
rect 22090 22820 22094 22876
rect 22030 22816 22094 22820
rect 28736 22876 28800 22880
rect 28736 22820 28740 22876
rect 28740 22820 28796 22876
rect 28796 22820 28800 22876
rect 28736 22816 28800 22820
rect 28816 22876 28880 22880
rect 28816 22820 28820 22876
rect 28820 22820 28876 22876
rect 28876 22820 28880 22876
rect 28816 22816 28880 22820
rect 28896 22876 28960 22880
rect 28896 22820 28900 22876
rect 28900 22820 28956 22876
rect 28956 22820 28960 22876
rect 28896 22816 28960 22820
rect 28976 22876 29040 22880
rect 28976 22820 28980 22876
rect 28980 22820 29036 22876
rect 29036 22820 29040 22876
rect 28976 22816 29040 22820
rect 4425 22332 4489 22336
rect 4425 22276 4429 22332
rect 4429 22276 4485 22332
rect 4485 22276 4489 22332
rect 4425 22272 4489 22276
rect 4505 22332 4569 22336
rect 4505 22276 4509 22332
rect 4509 22276 4565 22332
rect 4565 22276 4569 22332
rect 4505 22272 4569 22276
rect 4585 22332 4649 22336
rect 4585 22276 4589 22332
rect 4589 22276 4645 22332
rect 4645 22276 4649 22332
rect 4585 22272 4649 22276
rect 4665 22332 4729 22336
rect 4665 22276 4669 22332
rect 4669 22276 4725 22332
rect 4725 22276 4729 22332
rect 4665 22272 4729 22276
rect 11371 22332 11435 22336
rect 11371 22276 11375 22332
rect 11375 22276 11431 22332
rect 11431 22276 11435 22332
rect 11371 22272 11435 22276
rect 11451 22332 11515 22336
rect 11451 22276 11455 22332
rect 11455 22276 11511 22332
rect 11511 22276 11515 22332
rect 11451 22272 11515 22276
rect 11531 22332 11595 22336
rect 11531 22276 11535 22332
rect 11535 22276 11591 22332
rect 11591 22276 11595 22332
rect 11531 22272 11595 22276
rect 11611 22332 11675 22336
rect 11611 22276 11615 22332
rect 11615 22276 11671 22332
rect 11671 22276 11675 22332
rect 11611 22272 11675 22276
rect 18317 22332 18381 22336
rect 18317 22276 18321 22332
rect 18321 22276 18377 22332
rect 18377 22276 18381 22332
rect 18317 22272 18381 22276
rect 18397 22332 18461 22336
rect 18397 22276 18401 22332
rect 18401 22276 18457 22332
rect 18457 22276 18461 22332
rect 18397 22272 18461 22276
rect 18477 22332 18541 22336
rect 18477 22276 18481 22332
rect 18481 22276 18537 22332
rect 18537 22276 18541 22332
rect 18477 22272 18541 22276
rect 18557 22332 18621 22336
rect 18557 22276 18561 22332
rect 18561 22276 18617 22332
rect 18617 22276 18621 22332
rect 18557 22272 18621 22276
rect 25263 22332 25327 22336
rect 25263 22276 25267 22332
rect 25267 22276 25323 22332
rect 25323 22276 25327 22332
rect 25263 22272 25327 22276
rect 25343 22332 25407 22336
rect 25343 22276 25347 22332
rect 25347 22276 25403 22332
rect 25403 22276 25407 22332
rect 25343 22272 25407 22276
rect 25423 22332 25487 22336
rect 25423 22276 25427 22332
rect 25427 22276 25483 22332
rect 25483 22276 25487 22332
rect 25423 22272 25487 22276
rect 25503 22332 25567 22336
rect 25503 22276 25507 22332
rect 25507 22276 25563 22332
rect 25563 22276 25567 22332
rect 25503 22272 25567 22276
rect 7898 21788 7962 21792
rect 7898 21732 7902 21788
rect 7902 21732 7958 21788
rect 7958 21732 7962 21788
rect 7898 21728 7962 21732
rect 7978 21788 8042 21792
rect 7978 21732 7982 21788
rect 7982 21732 8038 21788
rect 8038 21732 8042 21788
rect 7978 21728 8042 21732
rect 8058 21788 8122 21792
rect 8058 21732 8062 21788
rect 8062 21732 8118 21788
rect 8118 21732 8122 21788
rect 8058 21728 8122 21732
rect 8138 21788 8202 21792
rect 8138 21732 8142 21788
rect 8142 21732 8198 21788
rect 8198 21732 8202 21788
rect 8138 21728 8202 21732
rect 14844 21788 14908 21792
rect 14844 21732 14848 21788
rect 14848 21732 14904 21788
rect 14904 21732 14908 21788
rect 14844 21728 14908 21732
rect 14924 21788 14988 21792
rect 14924 21732 14928 21788
rect 14928 21732 14984 21788
rect 14984 21732 14988 21788
rect 14924 21728 14988 21732
rect 15004 21788 15068 21792
rect 15004 21732 15008 21788
rect 15008 21732 15064 21788
rect 15064 21732 15068 21788
rect 15004 21728 15068 21732
rect 15084 21788 15148 21792
rect 15084 21732 15088 21788
rect 15088 21732 15144 21788
rect 15144 21732 15148 21788
rect 15084 21728 15148 21732
rect 21790 21788 21854 21792
rect 21790 21732 21794 21788
rect 21794 21732 21850 21788
rect 21850 21732 21854 21788
rect 21790 21728 21854 21732
rect 21870 21788 21934 21792
rect 21870 21732 21874 21788
rect 21874 21732 21930 21788
rect 21930 21732 21934 21788
rect 21870 21728 21934 21732
rect 21950 21788 22014 21792
rect 21950 21732 21954 21788
rect 21954 21732 22010 21788
rect 22010 21732 22014 21788
rect 21950 21728 22014 21732
rect 22030 21788 22094 21792
rect 22030 21732 22034 21788
rect 22034 21732 22090 21788
rect 22090 21732 22094 21788
rect 22030 21728 22094 21732
rect 28736 21788 28800 21792
rect 28736 21732 28740 21788
rect 28740 21732 28796 21788
rect 28796 21732 28800 21788
rect 28736 21728 28800 21732
rect 28816 21788 28880 21792
rect 28816 21732 28820 21788
rect 28820 21732 28876 21788
rect 28876 21732 28880 21788
rect 28816 21728 28880 21732
rect 28896 21788 28960 21792
rect 28896 21732 28900 21788
rect 28900 21732 28956 21788
rect 28956 21732 28960 21788
rect 28896 21728 28960 21732
rect 28976 21788 29040 21792
rect 28976 21732 28980 21788
rect 28980 21732 29036 21788
rect 29036 21732 29040 21788
rect 28976 21728 29040 21732
rect 4425 21244 4489 21248
rect 4425 21188 4429 21244
rect 4429 21188 4485 21244
rect 4485 21188 4489 21244
rect 4425 21184 4489 21188
rect 4505 21244 4569 21248
rect 4505 21188 4509 21244
rect 4509 21188 4565 21244
rect 4565 21188 4569 21244
rect 4505 21184 4569 21188
rect 4585 21244 4649 21248
rect 4585 21188 4589 21244
rect 4589 21188 4645 21244
rect 4645 21188 4649 21244
rect 4585 21184 4649 21188
rect 4665 21244 4729 21248
rect 4665 21188 4669 21244
rect 4669 21188 4725 21244
rect 4725 21188 4729 21244
rect 4665 21184 4729 21188
rect 11371 21244 11435 21248
rect 11371 21188 11375 21244
rect 11375 21188 11431 21244
rect 11431 21188 11435 21244
rect 11371 21184 11435 21188
rect 11451 21244 11515 21248
rect 11451 21188 11455 21244
rect 11455 21188 11511 21244
rect 11511 21188 11515 21244
rect 11451 21184 11515 21188
rect 11531 21244 11595 21248
rect 11531 21188 11535 21244
rect 11535 21188 11591 21244
rect 11591 21188 11595 21244
rect 11531 21184 11595 21188
rect 11611 21244 11675 21248
rect 11611 21188 11615 21244
rect 11615 21188 11671 21244
rect 11671 21188 11675 21244
rect 11611 21184 11675 21188
rect 18317 21244 18381 21248
rect 18317 21188 18321 21244
rect 18321 21188 18377 21244
rect 18377 21188 18381 21244
rect 18317 21184 18381 21188
rect 18397 21244 18461 21248
rect 18397 21188 18401 21244
rect 18401 21188 18457 21244
rect 18457 21188 18461 21244
rect 18397 21184 18461 21188
rect 18477 21244 18541 21248
rect 18477 21188 18481 21244
rect 18481 21188 18537 21244
rect 18537 21188 18541 21244
rect 18477 21184 18541 21188
rect 18557 21244 18621 21248
rect 18557 21188 18561 21244
rect 18561 21188 18617 21244
rect 18617 21188 18621 21244
rect 18557 21184 18621 21188
rect 25263 21244 25327 21248
rect 25263 21188 25267 21244
rect 25267 21188 25323 21244
rect 25323 21188 25327 21244
rect 25263 21184 25327 21188
rect 25343 21244 25407 21248
rect 25343 21188 25347 21244
rect 25347 21188 25403 21244
rect 25403 21188 25407 21244
rect 25343 21184 25407 21188
rect 25423 21244 25487 21248
rect 25423 21188 25427 21244
rect 25427 21188 25483 21244
rect 25483 21188 25487 21244
rect 25423 21184 25487 21188
rect 25503 21244 25567 21248
rect 25503 21188 25507 21244
rect 25507 21188 25563 21244
rect 25563 21188 25567 21244
rect 25503 21184 25567 21188
rect 7898 20700 7962 20704
rect 7898 20644 7902 20700
rect 7902 20644 7958 20700
rect 7958 20644 7962 20700
rect 7898 20640 7962 20644
rect 7978 20700 8042 20704
rect 7978 20644 7982 20700
rect 7982 20644 8038 20700
rect 8038 20644 8042 20700
rect 7978 20640 8042 20644
rect 8058 20700 8122 20704
rect 8058 20644 8062 20700
rect 8062 20644 8118 20700
rect 8118 20644 8122 20700
rect 8058 20640 8122 20644
rect 8138 20700 8202 20704
rect 8138 20644 8142 20700
rect 8142 20644 8198 20700
rect 8198 20644 8202 20700
rect 8138 20640 8202 20644
rect 14844 20700 14908 20704
rect 14844 20644 14848 20700
rect 14848 20644 14904 20700
rect 14904 20644 14908 20700
rect 14844 20640 14908 20644
rect 14924 20700 14988 20704
rect 14924 20644 14928 20700
rect 14928 20644 14984 20700
rect 14984 20644 14988 20700
rect 14924 20640 14988 20644
rect 15004 20700 15068 20704
rect 15004 20644 15008 20700
rect 15008 20644 15064 20700
rect 15064 20644 15068 20700
rect 15004 20640 15068 20644
rect 15084 20700 15148 20704
rect 15084 20644 15088 20700
rect 15088 20644 15144 20700
rect 15144 20644 15148 20700
rect 15084 20640 15148 20644
rect 21790 20700 21854 20704
rect 21790 20644 21794 20700
rect 21794 20644 21850 20700
rect 21850 20644 21854 20700
rect 21790 20640 21854 20644
rect 21870 20700 21934 20704
rect 21870 20644 21874 20700
rect 21874 20644 21930 20700
rect 21930 20644 21934 20700
rect 21870 20640 21934 20644
rect 21950 20700 22014 20704
rect 21950 20644 21954 20700
rect 21954 20644 22010 20700
rect 22010 20644 22014 20700
rect 21950 20640 22014 20644
rect 22030 20700 22094 20704
rect 22030 20644 22034 20700
rect 22034 20644 22090 20700
rect 22090 20644 22094 20700
rect 22030 20640 22094 20644
rect 28736 20700 28800 20704
rect 28736 20644 28740 20700
rect 28740 20644 28796 20700
rect 28796 20644 28800 20700
rect 28736 20640 28800 20644
rect 28816 20700 28880 20704
rect 28816 20644 28820 20700
rect 28820 20644 28876 20700
rect 28876 20644 28880 20700
rect 28816 20640 28880 20644
rect 28896 20700 28960 20704
rect 28896 20644 28900 20700
rect 28900 20644 28956 20700
rect 28956 20644 28960 20700
rect 28896 20640 28960 20644
rect 28976 20700 29040 20704
rect 28976 20644 28980 20700
rect 28980 20644 29036 20700
rect 29036 20644 29040 20700
rect 28976 20640 29040 20644
rect 4425 20156 4489 20160
rect 4425 20100 4429 20156
rect 4429 20100 4485 20156
rect 4485 20100 4489 20156
rect 4425 20096 4489 20100
rect 4505 20156 4569 20160
rect 4505 20100 4509 20156
rect 4509 20100 4565 20156
rect 4565 20100 4569 20156
rect 4505 20096 4569 20100
rect 4585 20156 4649 20160
rect 4585 20100 4589 20156
rect 4589 20100 4645 20156
rect 4645 20100 4649 20156
rect 4585 20096 4649 20100
rect 4665 20156 4729 20160
rect 4665 20100 4669 20156
rect 4669 20100 4725 20156
rect 4725 20100 4729 20156
rect 4665 20096 4729 20100
rect 11371 20156 11435 20160
rect 11371 20100 11375 20156
rect 11375 20100 11431 20156
rect 11431 20100 11435 20156
rect 11371 20096 11435 20100
rect 11451 20156 11515 20160
rect 11451 20100 11455 20156
rect 11455 20100 11511 20156
rect 11511 20100 11515 20156
rect 11451 20096 11515 20100
rect 11531 20156 11595 20160
rect 11531 20100 11535 20156
rect 11535 20100 11591 20156
rect 11591 20100 11595 20156
rect 11531 20096 11595 20100
rect 11611 20156 11675 20160
rect 11611 20100 11615 20156
rect 11615 20100 11671 20156
rect 11671 20100 11675 20156
rect 11611 20096 11675 20100
rect 18317 20156 18381 20160
rect 18317 20100 18321 20156
rect 18321 20100 18377 20156
rect 18377 20100 18381 20156
rect 18317 20096 18381 20100
rect 18397 20156 18461 20160
rect 18397 20100 18401 20156
rect 18401 20100 18457 20156
rect 18457 20100 18461 20156
rect 18397 20096 18461 20100
rect 18477 20156 18541 20160
rect 18477 20100 18481 20156
rect 18481 20100 18537 20156
rect 18537 20100 18541 20156
rect 18477 20096 18541 20100
rect 18557 20156 18621 20160
rect 18557 20100 18561 20156
rect 18561 20100 18617 20156
rect 18617 20100 18621 20156
rect 18557 20096 18621 20100
rect 25263 20156 25327 20160
rect 25263 20100 25267 20156
rect 25267 20100 25323 20156
rect 25323 20100 25327 20156
rect 25263 20096 25327 20100
rect 25343 20156 25407 20160
rect 25343 20100 25347 20156
rect 25347 20100 25403 20156
rect 25403 20100 25407 20156
rect 25343 20096 25407 20100
rect 25423 20156 25487 20160
rect 25423 20100 25427 20156
rect 25427 20100 25483 20156
rect 25483 20100 25487 20156
rect 25423 20096 25487 20100
rect 25503 20156 25567 20160
rect 25503 20100 25507 20156
rect 25507 20100 25563 20156
rect 25563 20100 25567 20156
rect 25503 20096 25567 20100
rect 7898 19612 7962 19616
rect 7898 19556 7902 19612
rect 7902 19556 7958 19612
rect 7958 19556 7962 19612
rect 7898 19552 7962 19556
rect 7978 19612 8042 19616
rect 7978 19556 7982 19612
rect 7982 19556 8038 19612
rect 8038 19556 8042 19612
rect 7978 19552 8042 19556
rect 8058 19612 8122 19616
rect 8058 19556 8062 19612
rect 8062 19556 8118 19612
rect 8118 19556 8122 19612
rect 8058 19552 8122 19556
rect 8138 19612 8202 19616
rect 8138 19556 8142 19612
rect 8142 19556 8198 19612
rect 8198 19556 8202 19612
rect 8138 19552 8202 19556
rect 14844 19612 14908 19616
rect 14844 19556 14848 19612
rect 14848 19556 14904 19612
rect 14904 19556 14908 19612
rect 14844 19552 14908 19556
rect 14924 19612 14988 19616
rect 14924 19556 14928 19612
rect 14928 19556 14984 19612
rect 14984 19556 14988 19612
rect 14924 19552 14988 19556
rect 15004 19612 15068 19616
rect 15004 19556 15008 19612
rect 15008 19556 15064 19612
rect 15064 19556 15068 19612
rect 15004 19552 15068 19556
rect 15084 19612 15148 19616
rect 15084 19556 15088 19612
rect 15088 19556 15144 19612
rect 15144 19556 15148 19612
rect 15084 19552 15148 19556
rect 21790 19612 21854 19616
rect 21790 19556 21794 19612
rect 21794 19556 21850 19612
rect 21850 19556 21854 19612
rect 21790 19552 21854 19556
rect 21870 19612 21934 19616
rect 21870 19556 21874 19612
rect 21874 19556 21930 19612
rect 21930 19556 21934 19612
rect 21870 19552 21934 19556
rect 21950 19612 22014 19616
rect 21950 19556 21954 19612
rect 21954 19556 22010 19612
rect 22010 19556 22014 19612
rect 21950 19552 22014 19556
rect 22030 19612 22094 19616
rect 22030 19556 22034 19612
rect 22034 19556 22090 19612
rect 22090 19556 22094 19612
rect 22030 19552 22094 19556
rect 28736 19612 28800 19616
rect 28736 19556 28740 19612
rect 28740 19556 28796 19612
rect 28796 19556 28800 19612
rect 28736 19552 28800 19556
rect 28816 19612 28880 19616
rect 28816 19556 28820 19612
rect 28820 19556 28876 19612
rect 28876 19556 28880 19612
rect 28816 19552 28880 19556
rect 28896 19612 28960 19616
rect 28896 19556 28900 19612
rect 28900 19556 28956 19612
rect 28956 19556 28960 19612
rect 28896 19552 28960 19556
rect 28976 19612 29040 19616
rect 28976 19556 28980 19612
rect 28980 19556 29036 19612
rect 29036 19556 29040 19612
rect 28976 19552 29040 19556
rect 4425 19068 4489 19072
rect 4425 19012 4429 19068
rect 4429 19012 4485 19068
rect 4485 19012 4489 19068
rect 4425 19008 4489 19012
rect 4505 19068 4569 19072
rect 4505 19012 4509 19068
rect 4509 19012 4565 19068
rect 4565 19012 4569 19068
rect 4505 19008 4569 19012
rect 4585 19068 4649 19072
rect 4585 19012 4589 19068
rect 4589 19012 4645 19068
rect 4645 19012 4649 19068
rect 4585 19008 4649 19012
rect 4665 19068 4729 19072
rect 4665 19012 4669 19068
rect 4669 19012 4725 19068
rect 4725 19012 4729 19068
rect 4665 19008 4729 19012
rect 11371 19068 11435 19072
rect 11371 19012 11375 19068
rect 11375 19012 11431 19068
rect 11431 19012 11435 19068
rect 11371 19008 11435 19012
rect 11451 19068 11515 19072
rect 11451 19012 11455 19068
rect 11455 19012 11511 19068
rect 11511 19012 11515 19068
rect 11451 19008 11515 19012
rect 11531 19068 11595 19072
rect 11531 19012 11535 19068
rect 11535 19012 11591 19068
rect 11591 19012 11595 19068
rect 11531 19008 11595 19012
rect 11611 19068 11675 19072
rect 11611 19012 11615 19068
rect 11615 19012 11671 19068
rect 11671 19012 11675 19068
rect 11611 19008 11675 19012
rect 18317 19068 18381 19072
rect 18317 19012 18321 19068
rect 18321 19012 18377 19068
rect 18377 19012 18381 19068
rect 18317 19008 18381 19012
rect 18397 19068 18461 19072
rect 18397 19012 18401 19068
rect 18401 19012 18457 19068
rect 18457 19012 18461 19068
rect 18397 19008 18461 19012
rect 18477 19068 18541 19072
rect 18477 19012 18481 19068
rect 18481 19012 18537 19068
rect 18537 19012 18541 19068
rect 18477 19008 18541 19012
rect 18557 19068 18621 19072
rect 18557 19012 18561 19068
rect 18561 19012 18617 19068
rect 18617 19012 18621 19068
rect 18557 19008 18621 19012
rect 25263 19068 25327 19072
rect 25263 19012 25267 19068
rect 25267 19012 25323 19068
rect 25323 19012 25327 19068
rect 25263 19008 25327 19012
rect 25343 19068 25407 19072
rect 25343 19012 25347 19068
rect 25347 19012 25403 19068
rect 25403 19012 25407 19068
rect 25343 19008 25407 19012
rect 25423 19068 25487 19072
rect 25423 19012 25427 19068
rect 25427 19012 25483 19068
rect 25483 19012 25487 19068
rect 25423 19008 25487 19012
rect 25503 19068 25567 19072
rect 25503 19012 25507 19068
rect 25507 19012 25563 19068
rect 25563 19012 25567 19068
rect 25503 19008 25567 19012
rect 7898 18524 7962 18528
rect 7898 18468 7902 18524
rect 7902 18468 7958 18524
rect 7958 18468 7962 18524
rect 7898 18464 7962 18468
rect 7978 18524 8042 18528
rect 7978 18468 7982 18524
rect 7982 18468 8038 18524
rect 8038 18468 8042 18524
rect 7978 18464 8042 18468
rect 8058 18524 8122 18528
rect 8058 18468 8062 18524
rect 8062 18468 8118 18524
rect 8118 18468 8122 18524
rect 8058 18464 8122 18468
rect 8138 18524 8202 18528
rect 8138 18468 8142 18524
rect 8142 18468 8198 18524
rect 8198 18468 8202 18524
rect 8138 18464 8202 18468
rect 14844 18524 14908 18528
rect 14844 18468 14848 18524
rect 14848 18468 14904 18524
rect 14904 18468 14908 18524
rect 14844 18464 14908 18468
rect 14924 18524 14988 18528
rect 14924 18468 14928 18524
rect 14928 18468 14984 18524
rect 14984 18468 14988 18524
rect 14924 18464 14988 18468
rect 15004 18524 15068 18528
rect 15004 18468 15008 18524
rect 15008 18468 15064 18524
rect 15064 18468 15068 18524
rect 15004 18464 15068 18468
rect 15084 18524 15148 18528
rect 15084 18468 15088 18524
rect 15088 18468 15144 18524
rect 15144 18468 15148 18524
rect 15084 18464 15148 18468
rect 21790 18524 21854 18528
rect 21790 18468 21794 18524
rect 21794 18468 21850 18524
rect 21850 18468 21854 18524
rect 21790 18464 21854 18468
rect 21870 18524 21934 18528
rect 21870 18468 21874 18524
rect 21874 18468 21930 18524
rect 21930 18468 21934 18524
rect 21870 18464 21934 18468
rect 21950 18524 22014 18528
rect 21950 18468 21954 18524
rect 21954 18468 22010 18524
rect 22010 18468 22014 18524
rect 21950 18464 22014 18468
rect 22030 18524 22094 18528
rect 22030 18468 22034 18524
rect 22034 18468 22090 18524
rect 22090 18468 22094 18524
rect 22030 18464 22094 18468
rect 28736 18524 28800 18528
rect 28736 18468 28740 18524
rect 28740 18468 28796 18524
rect 28796 18468 28800 18524
rect 28736 18464 28800 18468
rect 28816 18524 28880 18528
rect 28816 18468 28820 18524
rect 28820 18468 28876 18524
rect 28876 18468 28880 18524
rect 28816 18464 28880 18468
rect 28896 18524 28960 18528
rect 28896 18468 28900 18524
rect 28900 18468 28956 18524
rect 28956 18468 28960 18524
rect 28896 18464 28960 18468
rect 28976 18524 29040 18528
rect 28976 18468 28980 18524
rect 28980 18468 29036 18524
rect 29036 18468 29040 18524
rect 28976 18464 29040 18468
rect 4425 17980 4489 17984
rect 4425 17924 4429 17980
rect 4429 17924 4485 17980
rect 4485 17924 4489 17980
rect 4425 17920 4489 17924
rect 4505 17980 4569 17984
rect 4505 17924 4509 17980
rect 4509 17924 4565 17980
rect 4565 17924 4569 17980
rect 4505 17920 4569 17924
rect 4585 17980 4649 17984
rect 4585 17924 4589 17980
rect 4589 17924 4645 17980
rect 4645 17924 4649 17980
rect 4585 17920 4649 17924
rect 4665 17980 4729 17984
rect 4665 17924 4669 17980
rect 4669 17924 4725 17980
rect 4725 17924 4729 17980
rect 4665 17920 4729 17924
rect 11371 17980 11435 17984
rect 11371 17924 11375 17980
rect 11375 17924 11431 17980
rect 11431 17924 11435 17980
rect 11371 17920 11435 17924
rect 11451 17980 11515 17984
rect 11451 17924 11455 17980
rect 11455 17924 11511 17980
rect 11511 17924 11515 17980
rect 11451 17920 11515 17924
rect 11531 17980 11595 17984
rect 11531 17924 11535 17980
rect 11535 17924 11591 17980
rect 11591 17924 11595 17980
rect 11531 17920 11595 17924
rect 11611 17980 11675 17984
rect 11611 17924 11615 17980
rect 11615 17924 11671 17980
rect 11671 17924 11675 17980
rect 11611 17920 11675 17924
rect 18317 17980 18381 17984
rect 18317 17924 18321 17980
rect 18321 17924 18377 17980
rect 18377 17924 18381 17980
rect 18317 17920 18381 17924
rect 18397 17980 18461 17984
rect 18397 17924 18401 17980
rect 18401 17924 18457 17980
rect 18457 17924 18461 17980
rect 18397 17920 18461 17924
rect 18477 17980 18541 17984
rect 18477 17924 18481 17980
rect 18481 17924 18537 17980
rect 18537 17924 18541 17980
rect 18477 17920 18541 17924
rect 18557 17980 18621 17984
rect 18557 17924 18561 17980
rect 18561 17924 18617 17980
rect 18617 17924 18621 17980
rect 18557 17920 18621 17924
rect 25263 17980 25327 17984
rect 25263 17924 25267 17980
rect 25267 17924 25323 17980
rect 25323 17924 25327 17980
rect 25263 17920 25327 17924
rect 25343 17980 25407 17984
rect 25343 17924 25347 17980
rect 25347 17924 25403 17980
rect 25403 17924 25407 17980
rect 25343 17920 25407 17924
rect 25423 17980 25487 17984
rect 25423 17924 25427 17980
rect 25427 17924 25483 17980
rect 25483 17924 25487 17980
rect 25423 17920 25487 17924
rect 25503 17980 25567 17984
rect 25503 17924 25507 17980
rect 25507 17924 25563 17980
rect 25563 17924 25567 17980
rect 25503 17920 25567 17924
rect 7898 17436 7962 17440
rect 7898 17380 7902 17436
rect 7902 17380 7958 17436
rect 7958 17380 7962 17436
rect 7898 17376 7962 17380
rect 7978 17436 8042 17440
rect 7978 17380 7982 17436
rect 7982 17380 8038 17436
rect 8038 17380 8042 17436
rect 7978 17376 8042 17380
rect 8058 17436 8122 17440
rect 8058 17380 8062 17436
rect 8062 17380 8118 17436
rect 8118 17380 8122 17436
rect 8058 17376 8122 17380
rect 8138 17436 8202 17440
rect 8138 17380 8142 17436
rect 8142 17380 8198 17436
rect 8198 17380 8202 17436
rect 8138 17376 8202 17380
rect 14844 17436 14908 17440
rect 14844 17380 14848 17436
rect 14848 17380 14904 17436
rect 14904 17380 14908 17436
rect 14844 17376 14908 17380
rect 14924 17436 14988 17440
rect 14924 17380 14928 17436
rect 14928 17380 14984 17436
rect 14984 17380 14988 17436
rect 14924 17376 14988 17380
rect 15004 17436 15068 17440
rect 15004 17380 15008 17436
rect 15008 17380 15064 17436
rect 15064 17380 15068 17436
rect 15004 17376 15068 17380
rect 15084 17436 15148 17440
rect 15084 17380 15088 17436
rect 15088 17380 15144 17436
rect 15144 17380 15148 17436
rect 15084 17376 15148 17380
rect 21790 17436 21854 17440
rect 21790 17380 21794 17436
rect 21794 17380 21850 17436
rect 21850 17380 21854 17436
rect 21790 17376 21854 17380
rect 21870 17436 21934 17440
rect 21870 17380 21874 17436
rect 21874 17380 21930 17436
rect 21930 17380 21934 17436
rect 21870 17376 21934 17380
rect 21950 17436 22014 17440
rect 21950 17380 21954 17436
rect 21954 17380 22010 17436
rect 22010 17380 22014 17436
rect 21950 17376 22014 17380
rect 22030 17436 22094 17440
rect 22030 17380 22034 17436
rect 22034 17380 22090 17436
rect 22090 17380 22094 17436
rect 22030 17376 22094 17380
rect 28736 17436 28800 17440
rect 28736 17380 28740 17436
rect 28740 17380 28796 17436
rect 28796 17380 28800 17436
rect 28736 17376 28800 17380
rect 28816 17436 28880 17440
rect 28816 17380 28820 17436
rect 28820 17380 28876 17436
rect 28876 17380 28880 17436
rect 28816 17376 28880 17380
rect 28896 17436 28960 17440
rect 28896 17380 28900 17436
rect 28900 17380 28956 17436
rect 28956 17380 28960 17436
rect 28896 17376 28960 17380
rect 28976 17436 29040 17440
rect 28976 17380 28980 17436
rect 28980 17380 29036 17436
rect 29036 17380 29040 17436
rect 28976 17376 29040 17380
rect 4425 16892 4489 16896
rect 4425 16836 4429 16892
rect 4429 16836 4485 16892
rect 4485 16836 4489 16892
rect 4425 16832 4489 16836
rect 4505 16892 4569 16896
rect 4505 16836 4509 16892
rect 4509 16836 4565 16892
rect 4565 16836 4569 16892
rect 4505 16832 4569 16836
rect 4585 16892 4649 16896
rect 4585 16836 4589 16892
rect 4589 16836 4645 16892
rect 4645 16836 4649 16892
rect 4585 16832 4649 16836
rect 4665 16892 4729 16896
rect 4665 16836 4669 16892
rect 4669 16836 4725 16892
rect 4725 16836 4729 16892
rect 4665 16832 4729 16836
rect 11371 16892 11435 16896
rect 11371 16836 11375 16892
rect 11375 16836 11431 16892
rect 11431 16836 11435 16892
rect 11371 16832 11435 16836
rect 11451 16892 11515 16896
rect 11451 16836 11455 16892
rect 11455 16836 11511 16892
rect 11511 16836 11515 16892
rect 11451 16832 11515 16836
rect 11531 16892 11595 16896
rect 11531 16836 11535 16892
rect 11535 16836 11591 16892
rect 11591 16836 11595 16892
rect 11531 16832 11595 16836
rect 11611 16892 11675 16896
rect 11611 16836 11615 16892
rect 11615 16836 11671 16892
rect 11671 16836 11675 16892
rect 11611 16832 11675 16836
rect 18317 16892 18381 16896
rect 18317 16836 18321 16892
rect 18321 16836 18377 16892
rect 18377 16836 18381 16892
rect 18317 16832 18381 16836
rect 18397 16892 18461 16896
rect 18397 16836 18401 16892
rect 18401 16836 18457 16892
rect 18457 16836 18461 16892
rect 18397 16832 18461 16836
rect 18477 16892 18541 16896
rect 18477 16836 18481 16892
rect 18481 16836 18537 16892
rect 18537 16836 18541 16892
rect 18477 16832 18541 16836
rect 18557 16892 18621 16896
rect 18557 16836 18561 16892
rect 18561 16836 18617 16892
rect 18617 16836 18621 16892
rect 18557 16832 18621 16836
rect 25263 16892 25327 16896
rect 25263 16836 25267 16892
rect 25267 16836 25323 16892
rect 25323 16836 25327 16892
rect 25263 16832 25327 16836
rect 25343 16892 25407 16896
rect 25343 16836 25347 16892
rect 25347 16836 25403 16892
rect 25403 16836 25407 16892
rect 25343 16832 25407 16836
rect 25423 16892 25487 16896
rect 25423 16836 25427 16892
rect 25427 16836 25483 16892
rect 25483 16836 25487 16892
rect 25423 16832 25487 16836
rect 25503 16892 25567 16896
rect 25503 16836 25507 16892
rect 25507 16836 25563 16892
rect 25563 16836 25567 16892
rect 25503 16832 25567 16836
rect 7898 16348 7962 16352
rect 7898 16292 7902 16348
rect 7902 16292 7958 16348
rect 7958 16292 7962 16348
rect 7898 16288 7962 16292
rect 7978 16348 8042 16352
rect 7978 16292 7982 16348
rect 7982 16292 8038 16348
rect 8038 16292 8042 16348
rect 7978 16288 8042 16292
rect 8058 16348 8122 16352
rect 8058 16292 8062 16348
rect 8062 16292 8118 16348
rect 8118 16292 8122 16348
rect 8058 16288 8122 16292
rect 8138 16348 8202 16352
rect 8138 16292 8142 16348
rect 8142 16292 8198 16348
rect 8198 16292 8202 16348
rect 8138 16288 8202 16292
rect 14844 16348 14908 16352
rect 14844 16292 14848 16348
rect 14848 16292 14904 16348
rect 14904 16292 14908 16348
rect 14844 16288 14908 16292
rect 14924 16348 14988 16352
rect 14924 16292 14928 16348
rect 14928 16292 14984 16348
rect 14984 16292 14988 16348
rect 14924 16288 14988 16292
rect 15004 16348 15068 16352
rect 15004 16292 15008 16348
rect 15008 16292 15064 16348
rect 15064 16292 15068 16348
rect 15004 16288 15068 16292
rect 15084 16348 15148 16352
rect 15084 16292 15088 16348
rect 15088 16292 15144 16348
rect 15144 16292 15148 16348
rect 15084 16288 15148 16292
rect 21790 16348 21854 16352
rect 21790 16292 21794 16348
rect 21794 16292 21850 16348
rect 21850 16292 21854 16348
rect 21790 16288 21854 16292
rect 21870 16348 21934 16352
rect 21870 16292 21874 16348
rect 21874 16292 21930 16348
rect 21930 16292 21934 16348
rect 21870 16288 21934 16292
rect 21950 16348 22014 16352
rect 21950 16292 21954 16348
rect 21954 16292 22010 16348
rect 22010 16292 22014 16348
rect 21950 16288 22014 16292
rect 22030 16348 22094 16352
rect 22030 16292 22034 16348
rect 22034 16292 22090 16348
rect 22090 16292 22094 16348
rect 22030 16288 22094 16292
rect 28736 16348 28800 16352
rect 28736 16292 28740 16348
rect 28740 16292 28796 16348
rect 28796 16292 28800 16348
rect 28736 16288 28800 16292
rect 28816 16348 28880 16352
rect 28816 16292 28820 16348
rect 28820 16292 28876 16348
rect 28876 16292 28880 16348
rect 28816 16288 28880 16292
rect 28896 16348 28960 16352
rect 28896 16292 28900 16348
rect 28900 16292 28956 16348
rect 28956 16292 28960 16348
rect 28896 16288 28960 16292
rect 28976 16348 29040 16352
rect 28976 16292 28980 16348
rect 28980 16292 29036 16348
rect 29036 16292 29040 16348
rect 28976 16288 29040 16292
rect 4425 15804 4489 15808
rect 4425 15748 4429 15804
rect 4429 15748 4485 15804
rect 4485 15748 4489 15804
rect 4425 15744 4489 15748
rect 4505 15804 4569 15808
rect 4505 15748 4509 15804
rect 4509 15748 4565 15804
rect 4565 15748 4569 15804
rect 4505 15744 4569 15748
rect 4585 15804 4649 15808
rect 4585 15748 4589 15804
rect 4589 15748 4645 15804
rect 4645 15748 4649 15804
rect 4585 15744 4649 15748
rect 4665 15804 4729 15808
rect 4665 15748 4669 15804
rect 4669 15748 4725 15804
rect 4725 15748 4729 15804
rect 4665 15744 4729 15748
rect 11371 15804 11435 15808
rect 11371 15748 11375 15804
rect 11375 15748 11431 15804
rect 11431 15748 11435 15804
rect 11371 15744 11435 15748
rect 11451 15804 11515 15808
rect 11451 15748 11455 15804
rect 11455 15748 11511 15804
rect 11511 15748 11515 15804
rect 11451 15744 11515 15748
rect 11531 15804 11595 15808
rect 11531 15748 11535 15804
rect 11535 15748 11591 15804
rect 11591 15748 11595 15804
rect 11531 15744 11595 15748
rect 11611 15804 11675 15808
rect 11611 15748 11615 15804
rect 11615 15748 11671 15804
rect 11671 15748 11675 15804
rect 11611 15744 11675 15748
rect 18317 15804 18381 15808
rect 18317 15748 18321 15804
rect 18321 15748 18377 15804
rect 18377 15748 18381 15804
rect 18317 15744 18381 15748
rect 18397 15804 18461 15808
rect 18397 15748 18401 15804
rect 18401 15748 18457 15804
rect 18457 15748 18461 15804
rect 18397 15744 18461 15748
rect 18477 15804 18541 15808
rect 18477 15748 18481 15804
rect 18481 15748 18537 15804
rect 18537 15748 18541 15804
rect 18477 15744 18541 15748
rect 18557 15804 18621 15808
rect 18557 15748 18561 15804
rect 18561 15748 18617 15804
rect 18617 15748 18621 15804
rect 18557 15744 18621 15748
rect 25263 15804 25327 15808
rect 25263 15748 25267 15804
rect 25267 15748 25323 15804
rect 25323 15748 25327 15804
rect 25263 15744 25327 15748
rect 25343 15804 25407 15808
rect 25343 15748 25347 15804
rect 25347 15748 25403 15804
rect 25403 15748 25407 15804
rect 25343 15744 25407 15748
rect 25423 15804 25487 15808
rect 25423 15748 25427 15804
rect 25427 15748 25483 15804
rect 25483 15748 25487 15804
rect 25423 15744 25487 15748
rect 25503 15804 25567 15808
rect 25503 15748 25507 15804
rect 25507 15748 25563 15804
rect 25563 15748 25567 15804
rect 25503 15744 25567 15748
rect 7898 15260 7962 15264
rect 7898 15204 7902 15260
rect 7902 15204 7958 15260
rect 7958 15204 7962 15260
rect 7898 15200 7962 15204
rect 7978 15260 8042 15264
rect 7978 15204 7982 15260
rect 7982 15204 8038 15260
rect 8038 15204 8042 15260
rect 7978 15200 8042 15204
rect 8058 15260 8122 15264
rect 8058 15204 8062 15260
rect 8062 15204 8118 15260
rect 8118 15204 8122 15260
rect 8058 15200 8122 15204
rect 8138 15260 8202 15264
rect 8138 15204 8142 15260
rect 8142 15204 8198 15260
rect 8198 15204 8202 15260
rect 8138 15200 8202 15204
rect 14844 15260 14908 15264
rect 14844 15204 14848 15260
rect 14848 15204 14904 15260
rect 14904 15204 14908 15260
rect 14844 15200 14908 15204
rect 14924 15260 14988 15264
rect 14924 15204 14928 15260
rect 14928 15204 14984 15260
rect 14984 15204 14988 15260
rect 14924 15200 14988 15204
rect 15004 15260 15068 15264
rect 15004 15204 15008 15260
rect 15008 15204 15064 15260
rect 15064 15204 15068 15260
rect 15004 15200 15068 15204
rect 15084 15260 15148 15264
rect 15084 15204 15088 15260
rect 15088 15204 15144 15260
rect 15144 15204 15148 15260
rect 15084 15200 15148 15204
rect 21790 15260 21854 15264
rect 21790 15204 21794 15260
rect 21794 15204 21850 15260
rect 21850 15204 21854 15260
rect 21790 15200 21854 15204
rect 21870 15260 21934 15264
rect 21870 15204 21874 15260
rect 21874 15204 21930 15260
rect 21930 15204 21934 15260
rect 21870 15200 21934 15204
rect 21950 15260 22014 15264
rect 21950 15204 21954 15260
rect 21954 15204 22010 15260
rect 22010 15204 22014 15260
rect 21950 15200 22014 15204
rect 22030 15260 22094 15264
rect 22030 15204 22034 15260
rect 22034 15204 22090 15260
rect 22090 15204 22094 15260
rect 22030 15200 22094 15204
rect 28736 15260 28800 15264
rect 28736 15204 28740 15260
rect 28740 15204 28796 15260
rect 28796 15204 28800 15260
rect 28736 15200 28800 15204
rect 28816 15260 28880 15264
rect 28816 15204 28820 15260
rect 28820 15204 28876 15260
rect 28876 15204 28880 15260
rect 28816 15200 28880 15204
rect 28896 15260 28960 15264
rect 28896 15204 28900 15260
rect 28900 15204 28956 15260
rect 28956 15204 28960 15260
rect 28896 15200 28960 15204
rect 28976 15260 29040 15264
rect 28976 15204 28980 15260
rect 28980 15204 29036 15260
rect 29036 15204 29040 15260
rect 28976 15200 29040 15204
rect 4425 14716 4489 14720
rect 4425 14660 4429 14716
rect 4429 14660 4485 14716
rect 4485 14660 4489 14716
rect 4425 14656 4489 14660
rect 4505 14716 4569 14720
rect 4505 14660 4509 14716
rect 4509 14660 4565 14716
rect 4565 14660 4569 14716
rect 4505 14656 4569 14660
rect 4585 14716 4649 14720
rect 4585 14660 4589 14716
rect 4589 14660 4645 14716
rect 4645 14660 4649 14716
rect 4585 14656 4649 14660
rect 4665 14716 4729 14720
rect 4665 14660 4669 14716
rect 4669 14660 4725 14716
rect 4725 14660 4729 14716
rect 4665 14656 4729 14660
rect 11371 14716 11435 14720
rect 11371 14660 11375 14716
rect 11375 14660 11431 14716
rect 11431 14660 11435 14716
rect 11371 14656 11435 14660
rect 11451 14716 11515 14720
rect 11451 14660 11455 14716
rect 11455 14660 11511 14716
rect 11511 14660 11515 14716
rect 11451 14656 11515 14660
rect 11531 14716 11595 14720
rect 11531 14660 11535 14716
rect 11535 14660 11591 14716
rect 11591 14660 11595 14716
rect 11531 14656 11595 14660
rect 11611 14716 11675 14720
rect 11611 14660 11615 14716
rect 11615 14660 11671 14716
rect 11671 14660 11675 14716
rect 11611 14656 11675 14660
rect 18317 14716 18381 14720
rect 18317 14660 18321 14716
rect 18321 14660 18377 14716
rect 18377 14660 18381 14716
rect 18317 14656 18381 14660
rect 18397 14716 18461 14720
rect 18397 14660 18401 14716
rect 18401 14660 18457 14716
rect 18457 14660 18461 14716
rect 18397 14656 18461 14660
rect 18477 14716 18541 14720
rect 18477 14660 18481 14716
rect 18481 14660 18537 14716
rect 18537 14660 18541 14716
rect 18477 14656 18541 14660
rect 18557 14716 18621 14720
rect 18557 14660 18561 14716
rect 18561 14660 18617 14716
rect 18617 14660 18621 14716
rect 18557 14656 18621 14660
rect 25263 14716 25327 14720
rect 25263 14660 25267 14716
rect 25267 14660 25323 14716
rect 25323 14660 25327 14716
rect 25263 14656 25327 14660
rect 25343 14716 25407 14720
rect 25343 14660 25347 14716
rect 25347 14660 25403 14716
rect 25403 14660 25407 14716
rect 25343 14656 25407 14660
rect 25423 14716 25487 14720
rect 25423 14660 25427 14716
rect 25427 14660 25483 14716
rect 25483 14660 25487 14716
rect 25423 14656 25487 14660
rect 25503 14716 25567 14720
rect 25503 14660 25507 14716
rect 25507 14660 25563 14716
rect 25563 14660 25567 14716
rect 25503 14656 25567 14660
rect 7898 14172 7962 14176
rect 7898 14116 7902 14172
rect 7902 14116 7958 14172
rect 7958 14116 7962 14172
rect 7898 14112 7962 14116
rect 7978 14172 8042 14176
rect 7978 14116 7982 14172
rect 7982 14116 8038 14172
rect 8038 14116 8042 14172
rect 7978 14112 8042 14116
rect 8058 14172 8122 14176
rect 8058 14116 8062 14172
rect 8062 14116 8118 14172
rect 8118 14116 8122 14172
rect 8058 14112 8122 14116
rect 8138 14172 8202 14176
rect 8138 14116 8142 14172
rect 8142 14116 8198 14172
rect 8198 14116 8202 14172
rect 8138 14112 8202 14116
rect 14844 14172 14908 14176
rect 14844 14116 14848 14172
rect 14848 14116 14904 14172
rect 14904 14116 14908 14172
rect 14844 14112 14908 14116
rect 14924 14172 14988 14176
rect 14924 14116 14928 14172
rect 14928 14116 14984 14172
rect 14984 14116 14988 14172
rect 14924 14112 14988 14116
rect 15004 14172 15068 14176
rect 15004 14116 15008 14172
rect 15008 14116 15064 14172
rect 15064 14116 15068 14172
rect 15004 14112 15068 14116
rect 15084 14172 15148 14176
rect 15084 14116 15088 14172
rect 15088 14116 15144 14172
rect 15144 14116 15148 14172
rect 15084 14112 15148 14116
rect 21790 14172 21854 14176
rect 21790 14116 21794 14172
rect 21794 14116 21850 14172
rect 21850 14116 21854 14172
rect 21790 14112 21854 14116
rect 21870 14172 21934 14176
rect 21870 14116 21874 14172
rect 21874 14116 21930 14172
rect 21930 14116 21934 14172
rect 21870 14112 21934 14116
rect 21950 14172 22014 14176
rect 21950 14116 21954 14172
rect 21954 14116 22010 14172
rect 22010 14116 22014 14172
rect 21950 14112 22014 14116
rect 22030 14172 22094 14176
rect 22030 14116 22034 14172
rect 22034 14116 22090 14172
rect 22090 14116 22094 14172
rect 22030 14112 22094 14116
rect 28736 14172 28800 14176
rect 28736 14116 28740 14172
rect 28740 14116 28796 14172
rect 28796 14116 28800 14172
rect 28736 14112 28800 14116
rect 28816 14172 28880 14176
rect 28816 14116 28820 14172
rect 28820 14116 28876 14172
rect 28876 14116 28880 14172
rect 28816 14112 28880 14116
rect 28896 14172 28960 14176
rect 28896 14116 28900 14172
rect 28900 14116 28956 14172
rect 28956 14116 28960 14172
rect 28896 14112 28960 14116
rect 28976 14172 29040 14176
rect 28976 14116 28980 14172
rect 28980 14116 29036 14172
rect 29036 14116 29040 14172
rect 28976 14112 29040 14116
rect 4425 13628 4489 13632
rect 4425 13572 4429 13628
rect 4429 13572 4485 13628
rect 4485 13572 4489 13628
rect 4425 13568 4489 13572
rect 4505 13628 4569 13632
rect 4505 13572 4509 13628
rect 4509 13572 4565 13628
rect 4565 13572 4569 13628
rect 4505 13568 4569 13572
rect 4585 13628 4649 13632
rect 4585 13572 4589 13628
rect 4589 13572 4645 13628
rect 4645 13572 4649 13628
rect 4585 13568 4649 13572
rect 4665 13628 4729 13632
rect 4665 13572 4669 13628
rect 4669 13572 4725 13628
rect 4725 13572 4729 13628
rect 4665 13568 4729 13572
rect 11371 13628 11435 13632
rect 11371 13572 11375 13628
rect 11375 13572 11431 13628
rect 11431 13572 11435 13628
rect 11371 13568 11435 13572
rect 11451 13628 11515 13632
rect 11451 13572 11455 13628
rect 11455 13572 11511 13628
rect 11511 13572 11515 13628
rect 11451 13568 11515 13572
rect 11531 13628 11595 13632
rect 11531 13572 11535 13628
rect 11535 13572 11591 13628
rect 11591 13572 11595 13628
rect 11531 13568 11595 13572
rect 11611 13628 11675 13632
rect 11611 13572 11615 13628
rect 11615 13572 11671 13628
rect 11671 13572 11675 13628
rect 11611 13568 11675 13572
rect 18317 13628 18381 13632
rect 18317 13572 18321 13628
rect 18321 13572 18377 13628
rect 18377 13572 18381 13628
rect 18317 13568 18381 13572
rect 18397 13628 18461 13632
rect 18397 13572 18401 13628
rect 18401 13572 18457 13628
rect 18457 13572 18461 13628
rect 18397 13568 18461 13572
rect 18477 13628 18541 13632
rect 18477 13572 18481 13628
rect 18481 13572 18537 13628
rect 18537 13572 18541 13628
rect 18477 13568 18541 13572
rect 18557 13628 18621 13632
rect 18557 13572 18561 13628
rect 18561 13572 18617 13628
rect 18617 13572 18621 13628
rect 18557 13568 18621 13572
rect 25263 13628 25327 13632
rect 25263 13572 25267 13628
rect 25267 13572 25323 13628
rect 25323 13572 25327 13628
rect 25263 13568 25327 13572
rect 25343 13628 25407 13632
rect 25343 13572 25347 13628
rect 25347 13572 25403 13628
rect 25403 13572 25407 13628
rect 25343 13568 25407 13572
rect 25423 13628 25487 13632
rect 25423 13572 25427 13628
rect 25427 13572 25483 13628
rect 25483 13572 25487 13628
rect 25423 13568 25487 13572
rect 25503 13628 25567 13632
rect 25503 13572 25507 13628
rect 25507 13572 25563 13628
rect 25563 13572 25567 13628
rect 25503 13568 25567 13572
rect 7898 13084 7962 13088
rect 7898 13028 7902 13084
rect 7902 13028 7958 13084
rect 7958 13028 7962 13084
rect 7898 13024 7962 13028
rect 7978 13084 8042 13088
rect 7978 13028 7982 13084
rect 7982 13028 8038 13084
rect 8038 13028 8042 13084
rect 7978 13024 8042 13028
rect 8058 13084 8122 13088
rect 8058 13028 8062 13084
rect 8062 13028 8118 13084
rect 8118 13028 8122 13084
rect 8058 13024 8122 13028
rect 8138 13084 8202 13088
rect 8138 13028 8142 13084
rect 8142 13028 8198 13084
rect 8198 13028 8202 13084
rect 8138 13024 8202 13028
rect 14844 13084 14908 13088
rect 14844 13028 14848 13084
rect 14848 13028 14904 13084
rect 14904 13028 14908 13084
rect 14844 13024 14908 13028
rect 14924 13084 14988 13088
rect 14924 13028 14928 13084
rect 14928 13028 14984 13084
rect 14984 13028 14988 13084
rect 14924 13024 14988 13028
rect 15004 13084 15068 13088
rect 15004 13028 15008 13084
rect 15008 13028 15064 13084
rect 15064 13028 15068 13084
rect 15004 13024 15068 13028
rect 15084 13084 15148 13088
rect 15084 13028 15088 13084
rect 15088 13028 15144 13084
rect 15144 13028 15148 13084
rect 15084 13024 15148 13028
rect 21790 13084 21854 13088
rect 21790 13028 21794 13084
rect 21794 13028 21850 13084
rect 21850 13028 21854 13084
rect 21790 13024 21854 13028
rect 21870 13084 21934 13088
rect 21870 13028 21874 13084
rect 21874 13028 21930 13084
rect 21930 13028 21934 13084
rect 21870 13024 21934 13028
rect 21950 13084 22014 13088
rect 21950 13028 21954 13084
rect 21954 13028 22010 13084
rect 22010 13028 22014 13084
rect 21950 13024 22014 13028
rect 22030 13084 22094 13088
rect 22030 13028 22034 13084
rect 22034 13028 22090 13084
rect 22090 13028 22094 13084
rect 22030 13024 22094 13028
rect 28736 13084 28800 13088
rect 28736 13028 28740 13084
rect 28740 13028 28796 13084
rect 28796 13028 28800 13084
rect 28736 13024 28800 13028
rect 28816 13084 28880 13088
rect 28816 13028 28820 13084
rect 28820 13028 28876 13084
rect 28876 13028 28880 13084
rect 28816 13024 28880 13028
rect 28896 13084 28960 13088
rect 28896 13028 28900 13084
rect 28900 13028 28956 13084
rect 28956 13028 28960 13084
rect 28896 13024 28960 13028
rect 28976 13084 29040 13088
rect 28976 13028 28980 13084
rect 28980 13028 29036 13084
rect 29036 13028 29040 13084
rect 28976 13024 29040 13028
rect 4425 12540 4489 12544
rect 4425 12484 4429 12540
rect 4429 12484 4485 12540
rect 4485 12484 4489 12540
rect 4425 12480 4489 12484
rect 4505 12540 4569 12544
rect 4505 12484 4509 12540
rect 4509 12484 4565 12540
rect 4565 12484 4569 12540
rect 4505 12480 4569 12484
rect 4585 12540 4649 12544
rect 4585 12484 4589 12540
rect 4589 12484 4645 12540
rect 4645 12484 4649 12540
rect 4585 12480 4649 12484
rect 4665 12540 4729 12544
rect 4665 12484 4669 12540
rect 4669 12484 4725 12540
rect 4725 12484 4729 12540
rect 4665 12480 4729 12484
rect 11371 12540 11435 12544
rect 11371 12484 11375 12540
rect 11375 12484 11431 12540
rect 11431 12484 11435 12540
rect 11371 12480 11435 12484
rect 11451 12540 11515 12544
rect 11451 12484 11455 12540
rect 11455 12484 11511 12540
rect 11511 12484 11515 12540
rect 11451 12480 11515 12484
rect 11531 12540 11595 12544
rect 11531 12484 11535 12540
rect 11535 12484 11591 12540
rect 11591 12484 11595 12540
rect 11531 12480 11595 12484
rect 11611 12540 11675 12544
rect 11611 12484 11615 12540
rect 11615 12484 11671 12540
rect 11671 12484 11675 12540
rect 11611 12480 11675 12484
rect 18317 12540 18381 12544
rect 18317 12484 18321 12540
rect 18321 12484 18377 12540
rect 18377 12484 18381 12540
rect 18317 12480 18381 12484
rect 18397 12540 18461 12544
rect 18397 12484 18401 12540
rect 18401 12484 18457 12540
rect 18457 12484 18461 12540
rect 18397 12480 18461 12484
rect 18477 12540 18541 12544
rect 18477 12484 18481 12540
rect 18481 12484 18537 12540
rect 18537 12484 18541 12540
rect 18477 12480 18541 12484
rect 18557 12540 18621 12544
rect 18557 12484 18561 12540
rect 18561 12484 18617 12540
rect 18617 12484 18621 12540
rect 18557 12480 18621 12484
rect 25263 12540 25327 12544
rect 25263 12484 25267 12540
rect 25267 12484 25323 12540
rect 25323 12484 25327 12540
rect 25263 12480 25327 12484
rect 25343 12540 25407 12544
rect 25343 12484 25347 12540
rect 25347 12484 25403 12540
rect 25403 12484 25407 12540
rect 25343 12480 25407 12484
rect 25423 12540 25487 12544
rect 25423 12484 25427 12540
rect 25427 12484 25483 12540
rect 25483 12484 25487 12540
rect 25423 12480 25487 12484
rect 25503 12540 25567 12544
rect 25503 12484 25507 12540
rect 25507 12484 25563 12540
rect 25563 12484 25567 12540
rect 25503 12480 25567 12484
rect 7898 11996 7962 12000
rect 7898 11940 7902 11996
rect 7902 11940 7958 11996
rect 7958 11940 7962 11996
rect 7898 11936 7962 11940
rect 7978 11996 8042 12000
rect 7978 11940 7982 11996
rect 7982 11940 8038 11996
rect 8038 11940 8042 11996
rect 7978 11936 8042 11940
rect 8058 11996 8122 12000
rect 8058 11940 8062 11996
rect 8062 11940 8118 11996
rect 8118 11940 8122 11996
rect 8058 11936 8122 11940
rect 8138 11996 8202 12000
rect 8138 11940 8142 11996
rect 8142 11940 8198 11996
rect 8198 11940 8202 11996
rect 8138 11936 8202 11940
rect 14844 11996 14908 12000
rect 14844 11940 14848 11996
rect 14848 11940 14904 11996
rect 14904 11940 14908 11996
rect 14844 11936 14908 11940
rect 14924 11996 14988 12000
rect 14924 11940 14928 11996
rect 14928 11940 14984 11996
rect 14984 11940 14988 11996
rect 14924 11936 14988 11940
rect 15004 11996 15068 12000
rect 15004 11940 15008 11996
rect 15008 11940 15064 11996
rect 15064 11940 15068 11996
rect 15004 11936 15068 11940
rect 15084 11996 15148 12000
rect 15084 11940 15088 11996
rect 15088 11940 15144 11996
rect 15144 11940 15148 11996
rect 15084 11936 15148 11940
rect 21790 11996 21854 12000
rect 21790 11940 21794 11996
rect 21794 11940 21850 11996
rect 21850 11940 21854 11996
rect 21790 11936 21854 11940
rect 21870 11996 21934 12000
rect 21870 11940 21874 11996
rect 21874 11940 21930 11996
rect 21930 11940 21934 11996
rect 21870 11936 21934 11940
rect 21950 11996 22014 12000
rect 21950 11940 21954 11996
rect 21954 11940 22010 11996
rect 22010 11940 22014 11996
rect 21950 11936 22014 11940
rect 22030 11996 22094 12000
rect 22030 11940 22034 11996
rect 22034 11940 22090 11996
rect 22090 11940 22094 11996
rect 22030 11936 22094 11940
rect 28736 11996 28800 12000
rect 28736 11940 28740 11996
rect 28740 11940 28796 11996
rect 28796 11940 28800 11996
rect 28736 11936 28800 11940
rect 28816 11996 28880 12000
rect 28816 11940 28820 11996
rect 28820 11940 28876 11996
rect 28876 11940 28880 11996
rect 28816 11936 28880 11940
rect 28896 11996 28960 12000
rect 28896 11940 28900 11996
rect 28900 11940 28956 11996
rect 28956 11940 28960 11996
rect 28896 11936 28960 11940
rect 28976 11996 29040 12000
rect 28976 11940 28980 11996
rect 28980 11940 29036 11996
rect 29036 11940 29040 11996
rect 28976 11936 29040 11940
rect 4425 11452 4489 11456
rect 4425 11396 4429 11452
rect 4429 11396 4485 11452
rect 4485 11396 4489 11452
rect 4425 11392 4489 11396
rect 4505 11452 4569 11456
rect 4505 11396 4509 11452
rect 4509 11396 4565 11452
rect 4565 11396 4569 11452
rect 4505 11392 4569 11396
rect 4585 11452 4649 11456
rect 4585 11396 4589 11452
rect 4589 11396 4645 11452
rect 4645 11396 4649 11452
rect 4585 11392 4649 11396
rect 4665 11452 4729 11456
rect 4665 11396 4669 11452
rect 4669 11396 4725 11452
rect 4725 11396 4729 11452
rect 4665 11392 4729 11396
rect 11371 11452 11435 11456
rect 11371 11396 11375 11452
rect 11375 11396 11431 11452
rect 11431 11396 11435 11452
rect 11371 11392 11435 11396
rect 11451 11452 11515 11456
rect 11451 11396 11455 11452
rect 11455 11396 11511 11452
rect 11511 11396 11515 11452
rect 11451 11392 11515 11396
rect 11531 11452 11595 11456
rect 11531 11396 11535 11452
rect 11535 11396 11591 11452
rect 11591 11396 11595 11452
rect 11531 11392 11595 11396
rect 11611 11452 11675 11456
rect 11611 11396 11615 11452
rect 11615 11396 11671 11452
rect 11671 11396 11675 11452
rect 11611 11392 11675 11396
rect 18317 11452 18381 11456
rect 18317 11396 18321 11452
rect 18321 11396 18377 11452
rect 18377 11396 18381 11452
rect 18317 11392 18381 11396
rect 18397 11452 18461 11456
rect 18397 11396 18401 11452
rect 18401 11396 18457 11452
rect 18457 11396 18461 11452
rect 18397 11392 18461 11396
rect 18477 11452 18541 11456
rect 18477 11396 18481 11452
rect 18481 11396 18537 11452
rect 18537 11396 18541 11452
rect 18477 11392 18541 11396
rect 18557 11452 18621 11456
rect 18557 11396 18561 11452
rect 18561 11396 18617 11452
rect 18617 11396 18621 11452
rect 18557 11392 18621 11396
rect 25263 11452 25327 11456
rect 25263 11396 25267 11452
rect 25267 11396 25323 11452
rect 25323 11396 25327 11452
rect 25263 11392 25327 11396
rect 25343 11452 25407 11456
rect 25343 11396 25347 11452
rect 25347 11396 25403 11452
rect 25403 11396 25407 11452
rect 25343 11392 25407 11396
rect 25423 11452 25487 11456
rect 25423 11396 25427 11452
rect 25427 11396 25483 11452
rect 25483 11396 25487 11452
rect 25423 11392 25487 11396
rect 25503 11452 25567 11456
rect 25503 11396 25507 11452
rect 25507 11396 25563 11452
rect 25563 11396 25567 11452
rect 25503 11392 25567 11396
rect 7898 10908 7962 10912
rect 7898 10852 7902 10908
rect 7902 10852 7958 10908
rect 7958 10852 7962 10908
rect 7898 10848 7962 10852
rect 7978 10908 8042 10912
rect 7978 10852 7982 10908
rect 7982 10852 8038 10908
rect 8038 10852 8042 10908
rect 7978 10848 8042 10852
rect 8058 10908 8122 10912
rect 8058 10852 8062 10908
rect 8062 10852 8118 10908
rect 8118 10852 8122 10908
rect 8058 10848 8122 10852
rect 8138 10908 8202 10912
rect 8138 10852 8142 10908
rect 8142 10852 8198 10908
rect 8198 10852 8202 10908
rect 8138 10848 8202 10852
rect 14844 10908 14908 10912
rect 14844 10852 14848 10908
rect 14848 10852 14904 10908
rect 14904 10852 14908 10908
rect 14844 10848 14908 10852
rect 14924 10908 14988 10912
rect 14924 10852 14928 10908
rect 14928 10852 14984 10908
rect 14984 10852 14988 10908
rect 14924 10848 14988 10852
rect 15004 10908 15068 10912
rect 15004 10852 15008 10908
rect 15008 10852 15064 10908
rect 15064 10852 15068 10908
rect 15004 10848 15068 10852
rect 15084 10908 15148 10912
rect 15084 10852 15088 10908
rect 15088 10852 15144 10908
rect 15144 10852 15148 10908
rect 15084 10848 15148 10852
rect 21790 10908 21854 10912
rect 21790 10852 21794 10908
rect 21794 10852 21850 10908
rect 21850 10852 21854 10908
rect 21790 10848 21854 10852
rect 21870 10908 21934 10912
rect 21870 10852 21874 10908
rect 21874 10852 21930 10908
rect 21930 10852 21934 10908
rect 21870 10848 21934 10852
rect 21950 10908 22014 10912
rect 21950 10852 21954 10908
rect 21954 10852 22010 10908
rect 22010 10852 22014 10908
rect 21950 10848 22014 10852
rect 22030 10908 22094 10912
rect 22030 10852 22034 10908
rect 22034 10852 22090 10908
rect 22090 10852 22094 10908
rect 22030 10848 22094 10852
rect 28736 10908 28800 10912
rect 28736 10852 28740 10908
rect 28740 10852 28796 10908
rect 28796 10852 28800 10908
rect 28736 10848 28800 10852
rect 28816 10908 28880 10912
rect 28816 10852 28820 10908
rect 28820 10852 28876 10908
rect 28876 10852 28880 10908
rect 28816 10848 28880 10852
rect 28896 10908 28960 10912
rect 28896 10852 28900 10908
rect 28900 10852 28956 10908
rect 28956 10852 28960 10908
rect 28896 10848 28960 10852
rect 28976 10908 29040 10912
rect 28976 10852 28980 10908
rect 28980 10852 29036 10908
rect 29036 10852 29040 10908
rect 28976 10848 29040 10852
rect 4425 10364 4489 10368
rect 4425 10308 4429 10364
rect 4429 10308 4485 10364
rect 4485 10308 4489 10364
rect 4425 10304 4489 10308
rect 4505 10364 4569 10368
rect 4505 10308 4509 10364
rect 4509 10308 4565 10364
rect 4565 10308 4569 10364
rect 4505 10304 4569 10308
rect 4585 10364 4649 10368
rect 4585 10308 4589 10364
rect 4589 10308 4645 10364
rect 4645 10308 4649 10364
rect 4585 10304 4649 10308
rect 4665 10364 4729 10368
rect 4665 10308 4669 10364
rect 4669 10308 4725 10364
rect 4725 10308 4729 10364
rect 4665 10304 4729 10308
rect 11371 10364 11435 10368
rect 11371 10308 11375 10364
rect 11375 10308 11431 10364
rect 11431 10308 11435 10364
rect 11371 10304 11435 10308
rect 11451 10364 11515 10368
rect 11451 10308 11455 10364
rect 11455 10308 11511 10364
rect 11511 10308 11515 10364
rect 11451 10304 11515 10308
rect 11531 10364 11595 10368
rect 11531 10308 11535 10364
rect 11535 10308 11591 10364
rect 11591 10308 11595 10364
rect 11531 10304 11595 10308
rect 11611 10364 11675 10368
rect 11611 10308 11615 10364
rect 11615 10308 11671 10364
rect 11671 10308 11675 10364
rect 11611 10304 11675 10308
rect 18317 10364 18381 10368
rect 18317 10308 18321 10364
rect 18321 10308 18377 10364
rect 18377 10308 18381 10364
rect 18317 10304 18381 10308
rect 18397 10364 18461 10368
rect 18397 10308 18401 10364
rect 18401 10308 18457 10364
rect 18457 10308 18461 10364
rect 18397 10304 18461 10308
rect 18477 10364 18541 10368
rect 18477 10308 18481 10364
rect 18481 10308 18537 10364
rect 18537 10308 18541 10364
rect 18477 10304 18541 10308
rect 18557 10364 18621 10368
rect 18557 10308 18561 10364
rect 18561 10308 18617 10364
rect 18617 10308 18621 10364
rect 18557 10304 18621 10308
rect 25263 10364 25327 10368
rect 25263 10308 25267 10364
rect 25267 10308 25323 10364
rect 25323 10308 25327 10364
rect 25263 10304 25327 10308
rect 25343 10364 25407 10368
rect 25343 10308 25347 10364
rect 25347 10308 25403 10364
rect 25403 10308 25407 10364
rect 25343 10304 25407 10308
rect 25423 10364 25487 10368
rect 25423 10308 25427 10364
rect 25427 10308 25483 10364
rect 25483 10308 25487 10364
rect 25423 10304 25487 10308
rect 25503 10364 25567 10368
rect 25503 10308 25507 10364
rect 25507 10308 25563 10364
rect 25563 10308 25567 10364
rect 25503 10304 25567 10308
rect 7898 9820 7962 9824
rect 7898 9764 7902 9820
rect 7902 9764 7958 9820
rect 7958 9764 7962 9820
rect 7898 9760 7962 9764
rect 7978 9820 8042 9824
rect 7978 9764 7982 9820
rect 7982 9764 8038 9820
rect 8038 9764 8042 9820
rect 7978 9760 8042 9764
rect 8058 9820 8122 9824
rect 8058 9764 8062 9820
rect 8062 9764 8118 9820
rect 8118 9764 8122 9820
rect 8058 9760 8122 9764
rect 8138 9820 8202 9824
rect 8138 9764 8142 9820
rect 8142 9764 8198 9820
rect 8198 9764 8202 9820
rect 8138 9760 8202 9764
rect 14844 9820 14908 9824
rect 14844 9764 14848 9820
rect 14848 9764 14904 9820
rect 14904 9764 14908 9820
rect 14844 9760 14908 9764
rect 14924 9820 14988 9824
rect 14924 9764 14928 9820
rect 14928 9764 14984 9820
rect 14984 9764 14988 9820
rect 14924 9760 14988 9764
rect 15004 9820 15068 9824
rect 15004 9764 15008 9820
rect 15008 9764 15064 9820
rect 15064 9764 15068 9820
rect 15004 9760 15068 9764
rect 15084 9820 15148 9824
rect 15084 9764 15088 9820
rect 15088 9764 15144 9820
rect 15144 9764 15148 9820
rect 15084 9760 15148 9764
rect 21790 9820 21854 9824
rect 21790 9764 21794 9820
rect 21794 9764 21850 9820
rect 21850 9764 21854 9820
rect 21790 9760 21854 9764
rect 21870 9820 21934 9824
rect 21870 9764 21874 9820
rect 21874 9764 21930 9820
rect 21930 9764 21934 9820
rect 21870 9760 21934 9764
rect 21950 9820 22014 9824
rect 21950 9764 21954 9820
rect 21954 9764 22010 9820
rect 22010 9764 22014 9820
rect 21950 9760 22014 9764
rect 22030 9820 22094 9824
rect 22030 9764 22034 9820
rect 22034 9764 22090 9820
rect 22090 9764 22094 9820
rect 22030 9760 22094 9764
rect 28736 9820 28800 9824
rect 28736 9764 28740 9820
rect 28740 9764 28796 9820
rect 28796 9764 28800 9820
rect 28736 9760 28800 9764
rect 28816 9820 28880 9824
rect 28816 9764 28820 9820
rect 28820 9764 28876 9820
rect 28876 9764 28880 9820
rect 28816 9760 28880 9764
rect 28896 9820 28960 9824
rect 28896 9764 28900 9820
rect 28900 9764 28956 9820
rect 28956 9764 28960 9820
rect 28896 9760 28960 9764
rect 28976 9820 29040 9824
rect 28976 9764 28980 9820
rect 28980 9764 29036 9820
rect 29036 9764 29040 9820
rect 28976 9760 29040 9764
rect 4425 9276 4489 9280
rect 4425 9220 4429 9276
rect 4429 9220 4485 9276
rect 4485 9220 4489 9276
rect 4425 9216 4489 9220
rect 4505 9276 4569 9280
rect 4505 9220 4509 9276
rect 4509 9220 4565 9276
rect 4565 9220 4569 9276
rect 4505 9216 4569 9220
rect 4585 9276 4649 9280
rect 4585 9220 4589 9276
rect 4589 9220 4645 9276
rect 4645 9220 4649 9276
rect 4585 9216 4649 9220
rect 4665 9276 4729 9280
rect 4665 9220 4669 9276
rect 4669 9220 4725 9276
rect 4725 9220 4729 9276
rect 4665 9216 4729 9220
rect 11371 9276 11435 9280
rect 11371 9220 11375 9276
rect 11375 9220 11431 9276
rect 11431 9220 11435 9276
rect 11371 9216 11435 9220
rect 11451 9276 11515 9280
rect 11451 9220 11455 9276
rect 11455 9220 11511 9276
rect 11511 9220 11515 9276
rect 11451 9216 11515 9220
rect 11531 9276 11595 9280
rect 11531 9220 11535 9276
rect 11535 9220 11591 9276
rect 11591 9220 11595 9276
rect 11531 9216 11595 9220
rect 11611 9276 11675 9280
rect 11611 9220 11615 9276
rect 11615 9220 11671 9276
rect 11671 9220 11675 9276
rect 11611 9216 11675 9220
rect 18317 9276 18381 9280
rect 18317 9220 18321 9276
rect 18321 9220 18377 9276
rect 18377 9220 18381 9276
rect 18317 9216 18381 9220
rect 18397 9276 18461 9280
rect 18397 9220 18401 9276
rect 18401 9220 18457 9276
rect 18457 9220 18461 9276
rect 18397 9216 18461 9220
rect 18477 9276 18541 9280
rect 18477 9220 18481 9276
rect 18481 9220 18537 9276
rect 18537 9220 18541 9276
rect 18477 9216 18541 9220
rect 18557 9276 18621 9280
rect 18557 9220 18561 9276
rect 18561 9220 18617 9276
rect 18617 9220 18621 9276
rect 18557 9216 18621 9220
rect 25263 9276 25327 9280
rect 25263 9220 25267 9276
rect 25267 9220 25323 9276
rect 25323 9220 25327 9276
rect 25263 9216 25327 9220
rect 25343 9276 25407 9280
rect 25343 9220 25347 9276
rect 25347 9220 25403 9276
rect 25403 9220 25407 9276
rect 25343 9216 25407 9220
rect 25423 9276 25487 9280
rect 25423 9220 25427 9276
rect 25427 9220 25483 9276
rect 25483 9220 25487 9276
rect 25423 9216 25487 9220
rect 25503 9276 25567 9280
rect 25503 9220 25507 9276
rect 25507 9220 25563 9276
rect 25563 9220 25567 9276
rect 25503 9216 25567 9220
rect 7898 8732 7962 8736
rect 7898 8676 7902 8732
rect 7902 8676 7958 8732
rect 7958 8676 7962 8732
rect 7898 8672 7962 8676
rect 7978 8732 8042 8736
rect 7978 8676 7982 8732
rect 7982 8676 8038 8732
rect 8038 8676 8042 8732
rect 7978 8672 8042 8676
rect 8058 8732 8122 8736
rect 8058 8676 8062 8732
rect 8062 8676 8118 8732
rect 8118 8676 8122 8732
rect 8058 8672 8122 8676
rect 8138 8732 8202 8736
rect 8138 8676 8142 8732
rect 8142 8676 8198 8732
rect 8198 8676 8202 8732
rect 8138 8672 8202 8676
rect 14844 8732 14908 8736
rect 14844 8676 14848 8732
rect 14848 8676 14904 8732
rect 14904 8676 14908 8732
rect 14844 8672 14908 8676
rect 14924 8732 14988 8736
rect 14924 8676 14928 8732
rect 14928 8676 14984 8732
rect 14984 8676 14988 8732
rect 14924 8672 14988 8676
rect 15004 8732 15068 8736
rect 15004 8676 15008 8732
rect 15008 8676 15064 8732
rect 15064 8676 15068 8732
rect 15004 8672 15068 8676
rect 15084 8732 15148 8736
rect 15084 8676 15088 8732
rect 15088 8676 15144 8732
rect 15144 8676 15148 8732
rect 15084 8672 15148 8676
rect 21790 8732 21854 8736
rect 21790 8676 21794 8732
rect 21794 8676 21850 8732
rect 21850 8676 21854 8732
rect 21790 8672 21854 8676
rect 21870 8732 21934 8736
rect 21870 8676 21874 8732
rect 21874 8676 21930 8732
rect 21930 8676 21934 8732
rect 21870 8672 21934 8676
rect 21950 8732 22014 8736
rect 21950 8676 21954 8732
rect 21954 8676 22010 8732
rect 22010 8676 22014 8732
rect 21950 8672 22014 8676
rect 22030 8732 22094 8736
rect 22030 8676 22034 8732
rect 22034 8676 22090 8732
rect 22090 8676 22094 8732
rect 22030 8672 22094 8676
rect 28736 8732 28800 8736
rect 28736 8676 28740 8732
rect 28740 8676 28796 8732
rect 28796 8676 28800 8732
rect 28736 8672 28800 8676
rect 28816 8732 28880 8736
rect 28816 8676 28820 8732
rect 28820 8676 28876 8732
rect 28876 8676 28880 8732
rect 28816 8672 28880 8676
rect 28896 8732 28960 8736
rect 28896 8676 28900 8732
rect 28900 8676 28956 8732
rect 28956 8676 28960 8732
rect 28896 8672 28960 8676
rect 28976 8732 29040 8736
rect 28976 8676 28980 8732
rect 28980 8676 29036 8732
rect 29036 8676 29040 8732
rect 28976 8672 29040 8676
rect 4425 8188 4489 8192
rect 4425 8132 4429 8188
rect 4429 8132 4485 8188
rect 4485 8132 4489 8188
rect 4425 8128 4489 8132
rect 4505 8188 4569 8192
rect 4505 8132 4509 8188
rect 4509 8132 4565 8188
rect 4565 8132 4569 8188
rect 4505 8128 4569 8132
rect 4585 8188 4649 8192
rect 4585 8132 4589 8188
rect 4589 8132 4645 8188
rect 4645 8132 4649 8188
rect 4585 8128 4649 8132
rect 4665 8188 4729 8192
rect 4665 8132 4669 8188
rect 4669 8132 4725 8188
rect 4725 8132 4729 8188
rect 4665 8128 4729 8132
rect 11371 8188 11435 8192
rect 11371 8132 11375 8188
rect 11375 8132 11431 8188
rect 11431 8132 11435 8188
rect 11371 8128 11435 8132
rect 11451 8188 11515 8192
rect 11451 8132 11455 8188
rect 11455 8132 11511 8188
rect 11511 8132 11515 8188
rect 11451 8128 11515 8132
rect 11531 8188 11595 8192
rect 11531 8132 11535 8188
rect 11535 8132 11591 8188
rect 11591 8132 11595 8188
rect 11531 8128 11595 8132
rect 11611 8188 11675 8192
rect 11611 8132 11615 8188
rect 11615 8132 11671 8188
rect 11671 8132 11675 8188
rect 11611 8128 11675 8132
rect 18317 8188 18381 8192
rect 18317 8132 18321 8188
rect 18321 8132 18377 8188
rect 18377 8132 18381 8188
rect 18317 8128 18381 8132
rect 18397 8188 18461 8192
rect 18397 8132 18401 8188
rect 18401 8132 18457 8188
rect 18457 8132 18461 8188
rect 18397 8128 18461 8132
rect 18477 8188 18541 8192
rect 18477 8132 18481 8188
rect 18481 8132 18537 8188
rect 18537 8132 18541 8188
rect 18477 8128 18541 8132
rect 18557 8188 18621 8192
rect 18557 8132 18561 8188
rect 18561 8132 18617 8188
rect 18617 8132 18621 8188
rect 18557 8128 18621 8132
rect 25263 8188 25327 8192
rect 25263 8132 25267 8188
rect 25267 8132 25323 8188
rect 25323 8132 25327 8188
rect 25263 8128 25327 8132
rect 25343 8188 25407 8192
rect 25343 8132 25347 8188
rect 25347 8132 25403 8188
rect 25403 8132 25407 8188
rect 25343 8128 25407 8132
rect 25423 8188 25487 8192
rect 25423 8132 25427 8188
rect 25427 8132 25483 8188
rect 25483 8132 25487 8188
rect 25423 8128 25487 8132
rect 25503 8188 25567 8192
rect 25503 8132 25507 8188
rect 25507 8132 25563 8188
rect 25563 8132 25567 8188
rect 25503 8128 25567 8132
rect 7898 7644 7962 7648
rect 7898 7588 7902 7644
rect 7902 7588 7958 7644
rect 7958 7588 7962 7644
rect 7898 7584 7962 7588
rect 7978 7644 8042 7648
rect 7978 7588 7982 7644
rect 7982 7588 8038 7644
rect 8038 7588 8042 7644
rect 7978 7584 8042 7588
rect 8058 7644 8122 7648
rect 8058 7588 8062 7644
rect 8062 7588 8118 7644
rect 8118 7588 8122 7644
rect 8058 7584 8122 7588
rect 8138 7644 8202 7648
rect 8138 7588 8142 7644
rect 8142 7588 8198 7644
rect 8198 7588 8202 7644
rect 8138 7584 8202 7588
rect 14844 7644 14908 7648
rect 14844 7588 14848 7644
rect 14848 7588 14904 7644
rect 14904 7588 14908 7644
rect 14844 7584 14908 7588
rect 14924 7644 14988 7648
rect 14924 7588 14928 7644
rect 14928 7588 14984 7644
rect 14984 7588 14988 7644
rect 14924 7584 14988 7588
rect 15004 7644 15068 7648
rect 15004 7588 15008 7644
rect 15008 7588 15064 7644
rect 15064 7588 15068 7644
rect 15004 7584 15068 7588
rect 15084 7644 15148 7648
rect 15084 7588 15088 7644
rect 15088 7588 15144 7644
rect 15144 7588 15148 7644
rect 15084 7584 15148 7588
rect 21790 7644 21854 7648
rect 21790 7588 21794 7644
rect 21794 7588 21850 7644
rect 21850 7588 21854 7644
rect 21790 7584 21854 7588
rect 21870 7644 21934 7648
rect 21870 7588 21874 7644
rect 21874 7588 21930 7644
rect 21930 7588 21934 7644
rect 21870 7584 21934 7588
rect 21950 7644 22014 7648
rect 21950 7588 21954 7644
rect 21954 7588 22010 7644
rect 22010 7588 22014 7644
rect 21950 7584 22014 7588
rect 22030 7644 22094 7648
rect 22030 7588 22034 7644
rect 22034 7588 22090 7644
rect 22090 7588 22094 7644
rect 22030 7584 22094 7588
rect 28736 7644 28800 7648
rect 28736 7588 28740 7644
rect 28740 7588 28796 7644
rect 28796 7588 28800 7644
rect 28736 7584 28800 7588
rect 28816 7644 28880 7648
rect 28816 7588 28820 7644
rect 28820 7588 28876 7644
rect 28876 7588 28880 7644
rect 28816 7584 28880 7588
rect 28896 7644 28960 7648
rect 28896 7588 28900 7644
rect 28900 7588 28956 7644
rect 28956 7588 28960 7644
rect 28896 7584 28960 7588
rect 28976 7644 29040 7648
rect 28976 7588 28980 7644
rect 28980 7588 29036 7644
rect 29036 7588 29040 7644
rect 28976 7584 29040 7588
rect 4425 7100 4489 7104
rect 4425 7044 4429 7100
rect 4429 7044 4485 7100
rect 4485 7044 4489 7100
rect 4425 7040 4489 7044
rect 4505 7100 4569 7104
rect 4505 7044 4509 7100
rect 4509 7044 4565 7100
rect 4565 7044 4569 7100
rect 4505 7040 4569 7044
rect 4585 7100 4649 7104
rect 4585 7044 4589 7100
rect 4589 7044 4645 7100
rect 4645 7044 4649 7100
rect 4585 7040 4649 7044
rect 4665 7100 4729 7104
rect 4665 7044 4669 7100
rect 4669 7044 4725 7100
rect 4725 7044 4729 7100
rect 4665 7040 4729 7044
rect 11371 7100 11435 7104
rect 11371 7044 11375 7100
rect 11375 7044 11431 7100
rect 11431 7044 11435 7100
rect 11371 7040 11435 7044
rect 11451 7100 11515 7104
rect 11451 7044 11455 7100
rect 11455 7044 11511 7100
rect 11511 7044 11515 7100
rect 11451 7040 11515 7044
rect 11531 7100 11595 7104
rect 11531 7044 11535 7100
rect 11535 7044 11591 7100
rect 11591 7044 11595 7100
rect 11531 7040 11595 7044
rect 11611 7100 11675 7104
rect 11611 7044 11615 7100
rect 11615 7044 11671 7100
rect 11671 7044 11675 7100
rect 11611 7040 11675 7044
rect 18317 7100 18381 7104
rect 18317 7044 18321 7100
rect 18321 7044 18377 7100
rect 18377 7044 18381 7100
rect 18317 7040 18381 7044
rect 18397 7100 18461 7104
rect 18397 7044 18401 7100
rect 18401 7044 18457 7100
rect 18457 7044 18461 7100
rect 18397 7040 18461 7044
rect 18477 7100 18541 7104
rect 18477 7044 18481 7100
rect 18481 7044 18537 7100
rect 18537 7044 18541 7100
rect 18477 7040 18541 7044
rect 18557 7100 18621 7104
rect 18557 7044 18561 7100
rect 18561 7044 18617 7100
rect 18617 7044 18621 7100
rect 18557 7040 18621 7044
rect 25263 7100 25327 7104
rect 25263 7044 25267 7100
rect 25267 7044 25323 7100
rect 25323 7044 25327 7100
rect 25263 7040 25327 7044
rect 25343 7100 25407 7104
rect 25343 7044 25347 7100
rect 25347 7044 25403 7100
rect 25403 7044 25407 7100
rect 25343 7040 25407 7044
rect 25423 7100 25487 7104
rect 25423 7044 25427 7100
rect 25427 7044 25483 7100
rect 25483 7044 25487 7100
rect 25423 7040 25487 7044
rect 25503 7100 25567 7104
rect 25503 7044 25507 7100
rect 25507 7044 25563 7100
rect 25563 7044 25567 7100
rect 25503 7040 25567 7044
rect 7898 6556 7962 6560
rect 7898 6500 7902 6556
rect 7902 6500 7958 6556
rect 7958 6500 7962 6556
rect 7898 6496 7962 6500
rect 7978 6556 8042 6560
rect 7978 6500 7982 6556
rect 7982 6500 8038 6556
rect 8038 6500 8042 6556
rect 7978 6496 8042 6500
rect 8058 6556 8122 6560
rect 8058 6500 8062 6556
rect 8062 6500 8118 6556
rect 8118 6500 8122 6556
rect 8058 6496 8122 6500
rect 8138 6556 8202 6560
rect 8138 6500 8142 6556
rect 8142 6500 8198 6556
rect 8198 6500 8202 6556
rect 8138 6496 8202 6500
rect 14844 6556 14908 6560
rect 14844 6500 14848 6556
rect 14848 6500 14904 6556
rect 14904 6500 14908 6556
rect 14844 6496 14908 6500
rect 14924 6556 14988 6560
rect 14924 6500 14928 6556
rect 14928 6500 14984 6556
rect 14984 6500 14988 6556
rect 14924 6496 14988 6500
rect 15004 6556 15068 6560
rect 15004 6500 15008 6556
rect 15008 6500 15064 6556
rect 15064 6500 15068 6556
rect 15004 6496 15068 6500
rect 15084 6556 15148 6560
rect 15084 6500 15088 6556
rect 15088 6500 15144 6556
rect 15144 6500 15148 6556
rect 15084 6496 15148 6500
rect 21790 6556 21854 6560
rect 21790 6500 21794 6556
rect 21794 6500 21850 6556
rect 21850 6500 21854 6556
rect 21790 6496 21854 6500
rect 21870 6556 21934 6560
rect 21870 6500 21874 6556
rect 21874 6500 21930 6556
rect 21930 6500 21934 6556
rect 21870 6496 21934 6500
rect 21950 6556 22014 6560
rect 21950 6500 21954 6556
rect 21954 6500 22010 6556
rect 22010 6500 22014 6556
rect 21950 6496 22014 6500
rect 22030 6556 22094 6560
rect 22030 6500 22034 6556
rect 22034 6500 22090 6556
rect 22090 6500 22094 6556
rect 22030 6496 22094 6500
rect 28736 6556 28800 6560
rect 28736 6500 28740 6556
rect 28740 6500 28796 6556
rect 28796 6500 28800 6556
rect 28736 6496 28800 6500
rect 28816 6556 28880 6560
rect 28816 6500 28820 6556
rect 28820 6500 28876 6556
rect 28876 6500 28880 6556
rect 28816 6496 28880 6500
rect 28896 6556 28960 6560
rect 28896 6500 28900 6556
rect 28900 6500 28956 6556
rect 28956 6500 28960 6556
rect 28896 6496 28960 6500
rect 28976 6556 29040 6560
rect 28976 6500 28980 6556
rect 28980 6500 29036 6556
rect 29036 6500 29040 6556
rect 28976 6496 29040 6500
rect 4425 6012 4489 6016
rect 4425 5956 4429 6012
rect 4429 5956 4485 6012
rect 4485 5956 4489 6012
rect 4425 5952 4489 5956
rect 4505 6012 4569 6016
rect 4505 5956 4509 6012
rect 4509 5956 4565 6012
rect 4565 5956 4569 6012
rect 4505 5952 4569 5956
rect 4585 6012 4649 6016
rect 4585 5956 4589 6012
rect 4589 5956 4645 6012
rect 4645 5956 4649 6012
rect 4585 5952 4649 5956
rect 4665 6012 4729 6016
rect 4665 5956 4669 6012
rect 4669 5956 4725 6012
rect 4725 5956 4729 6012
rect 4665 5952 4729 5956
rect 11371 6012 11435 6016
rect 11371 5956 11375 6012
rect 11375 5956 11431 6012
rect 11431 5956 11435 6012
rect 11371 5952 11435 5956
rect 11451 6012 11515 6016
rect 11451 5956 11455 6012
rect 11455 5956 11511 6012
rect 11511 5956 11515 6012
rect 11451 5952 11515 5956
rect 11531 6012 11595 6016
rect 11531 5956 11535 6012
rect 11535 5956 11591 6012
rect 11591 5956 11595 6012
rect 11531 5952 11595 5956
rect 11611 6012 11675 6016
rect 11611 5956 11615 6012
rect 11615 5956 11671 6012
rect 11671 5956 11675 6012
rect 11611 5952 11675 5956
rect 18317 6012 18381 6016
rect 18317 5956 18321 6012
rect 18321 5956 18377 6012
rect 18377 5956 18381 6012
rect 18317 5952 18381 5956
rect 18397 6012 18461 6016
rect 18397 5956 18401 6012
rect 18401 5956 18457 6012
rect 18457 5956 18461 6012
rect 18397 5952 18461 5956
rect 18477 6012 18541 6016
rect 18477 5956 18481 6012
rect 18481 5956 18537 6012
rect 18537 5956 18541 6012
rect 18477 5952 18541 5956
rect 18557 6012 18621 6016
rect 18557 5956 18561 6012
rect 18561 5956 18617 6012
rect 18617 5956 18621 6012
rect 18557 5952 18621 5956
rect 25263 6012 25327 6016
rect 25263 5956 25267 6012
rect 25267 5956 25323 6012
rect 25323 5956 25327 6012
rect 25263 5952 25327 5956
rect 25343 6012 25407 6016
rect 25343 5956 25347 6012
rect 25347 5956 25403 6012
rect 25403 5956 25407 6012
rect 25343 5952 25407 5956
rect 25423 6012 25487 6016
rect 25423 5956 25427 6012
rect 25427 5956 25483 6012
rect 25483 5956 25487 6012
rect 25423 5952 25487 5956
rect 25503 6012 25567 6016
rect 25503 5956 25507 6012
rect 25507 5956 25563 6012
rect 25563 5956 25567 6012
rect 25503 5952 25567 5956
rect 7898 5468 7962 5472
rect 7898 5412 7902 5468
rect 7902 5412 7958 5468
rect 7958 5412 7962 5468
rect 7898 5408 7962 5412
rect 7978 5468 8042 5472
rect 7978 5412 7982 5468
rect 7982 5412 8038 5468
rect 8038 5412 8042 5468
rect 7978 5408 8042 5412
rect 8058 5468 8122 5472
rect 8058 5412 8062 5468
rect 8062 5412 8118 5468
rect 8118 5412 8122 5468
rect 8058 5408 8122 5412
rect 8138 5468 8202 5472
rect 8138 5412 8142 5468
rect 8142 5412 8198 5468
rect 8198 5412 8202 5468
rect 8138 5408 8202 5412
rect 14844 5468 14908 5472
rect 14844 5412 14848 5468
rect 14848 5412 14904 5468
rect 14904 5412 14908 5468
rect 14844 5408 14908 5412
rect 14924 5468 14988 5472
rect 14924 5412 14928 5468
rect 14928 5412 14984 5468
rect 14984 5412 14988 5468
rect 14924 5408 14988 5412
rect 15004 5468 15068 5472
rect 15004 5412 15008 5468
rect 15008 5412 15064 5468
rect 15064 5412 15068 5468
rect 15004 5408 15068 5412
rect 15084 5468 15148 5472
rect 15084 5412 15088 5468
rect 15088 5412 15144 5468
rect 15144 5412 15148 5468
rect 15084 5408 15148 5412
rect 21790 5468 21854 5472
rect 21790 5412 21794 5468
rect 21794 5412 21850 5468
rect 21850 5412 21854 5468
rect 21790 5408 21854 5412
rect 21870 5468 21934 5472
rect 21870 5412 21874 5468
rect 21874 5412 21930 5468
rect 21930 5412 21934 5468
rect 21870 5408 21934 5412
rect 21950 5468 22014 5472
rect 21950 5412 21954 5468
rect 21954 5412 22010 5468
rect 22010 5412 22014 5468
rect 21950 5408 22014 5412
rect 22030 5468 22094 5472
rect 22030 5412 22034 5468
rect 22034 5412 22090 5468
rect 22090 5412 22094 5468
rect 22030 5408 22094 5412
rect 28736 5468 28800 5472
rect 28736 5412 28740 5468
rect 28740 5412 28796 5468
rect 28796 5412 28800 5468
rect 28736 5408 28800 5412
rect 28816 5468 28880 5472
rect 28816 5412 28820 5468
rect 28820 5412 28876 5468
rect 28876 5412 28880 5468
rect 28816 5408 28880 5412
rect 28896 5468 28960 5472
rect 28896 5412 28900 5468
rect 28900 5412 28956 5468
rect 28956 5412 28960 5468
rect 28896 5408 28960 5412
rect 28976 5468 29040 5472
rect 28976 5412 28980 5468
rect 28980 5412 29036 5468
rect 29036 5412 29040 5468
rect 28976 5408 29040 5412
rect 4425 4924 4489 4928
rect 4425 4868 4429 4924
rect 4429 4868 4485 4924
rect 4485 4868 4489 4924
rect 4425 4864 4489 4868
rect 4505 4924 4569 4928
rect 4505 4868 4509 4924
rect 4509 4868 4565 4924
rect 4565 4868 4569 4924
rect 4505 4864 4569 4868
rect 4585 4924 4649 4928
rect 4585 4868 4589 4924
rect 4589 4868 4645 4924
rect 4645 4868 4649 4924
rect 4585 4864 4649 4868
rect 4665 4924 4729 4928
rect 4665 4868 4669 4924
rect 4669 4868 4725 4924
rect 4725 4868 4729 4924
rect 4665 4864 4729 4868
rect 11371 4924 11435 4928
rect 11371 4868 11375 4924
rect 11375 4868 11431 4924
rect 11431 4868 11435 4924
rect 11371 4864 11435 4868
rect 11451 4924 11515 4928
rect 11451 4868 11455 4924
rect 11455 4868 11511 4924
rect 11511 4868 11515 4924
rect 11451 4864 11515 4868
rect 11531 4924 11595 4928
rect 11531 4868 11535 4924
rect 11535 4868 11591 4924
rect 11591 4868 11595 4924
rect 11531 4864 11595 4868
rect 11611 4924 11675 4928
rect 11611 4868 11615 4924
rect 11615 4868 11671 4924
rect 11671 4868 11675 4924
rect 11611 4864 11675 4868
rect 18317 4924 18381 4928
rect 18317 4868 18321 4924
rect 18321 4868 18377 4924
rect 18377 4868 18381 4924
rect 18317 4864 18381 4868
rect 18397 4924 18461 4928
rect 18397 4868 18401 4924
rect 18401 4868 18457 4924
rect 18457 4868 18461 4924
rect 18397 4864 18461 4868
rect 18477 4924 18541 4928
rect 18477 4868 18481 4924
rect 18481 4868 18537 4924
rect 18537 4868 18541 4924
rect 18477 4864 18541 4868
rect 18557 4924 18621 4928
rect 18557 4868 18561 4924
rect 18561 4868 18617 4924
rect 18617 4868 18621 4924
rect 18557 4864 18621 4868
rect 25263 4924 25327 4928
rect 25263 4868 25267 4924
rect 25267 4868 25323 4924
rect 25323 4868 25327 4924
rect 25263 4864 25327 4868
rect 25343 4924 25407 4928
rect 25343 4868 25347 4924
rect 25347 4868 25403 4924
rect 25403 4868 25407 4924
rect 25343 4864 25407 4868
rect 25423 4924 25487 4928
rect 25423 4868 25427 4924
rect 25427 4868 25483 4924
rect 25483 4868 25487 4924
rect 25423 4864 25487 4868
rect 25503 4924 25567 4928
rect 25503 4868 25507 4924
rect 25507 4868 25563 4924
rect 25563 4868 25567 4924
rect 25503 4864 25567 4868
rect 7898 4380 7962 4384
rect 7898 4324 7902 4380
rect 7902 4324 7958 4380
rect 7958 4324 7962 4380
rect 7898 4320 7962 4324
rect 7978 4380 8042 4384
rect 7978 4324 7982 4380
rect 7982 4324 8038 4380
rect 8038 4324 8042 4380
rect 7978 4320 8042 4324
rect 8058 4380 8122 4384
rect 8058 4324 8062 4380
rect 8062 4324 8118 4380
rect 8118 4324 8122 4380
rect 8058 4320 8122 4324
rect 8138 4380 8202 4384
rect 8138 4324 8142 4380
rect 8142 4324 8198 4380
rect 8198 4324 8202 4380
rect 8138 4320 8202 4324
rect 14844 4380 14908 4384
rect 14844 4324 14848 4380
rect 14848 4324 14904 4380
rect 14904 4324 14908 4380
rect 14844 4320 14908 4324
rect 14924 4380 14988 4384
rect 14924 4324 14928 4380
rect 14928 4324 14984 4380
rect 14984 4324 14988 4380
rect 14924 4320 14988 4324
rect 15004 4380 15068 4384
rect 15004 4324 15008 4380
rect 15008 4324 15064 4380
rect 15064 4324 15068 4380
rect 15004 4320 15068 4324
rect 15084 4380 15148 4384
rect 15084 4324 15088 4380
rect 15088 4324 15144 4380
rect 15144 4324 15148 4380
rect 15084 4320 15148 4324
rect 21790 4380 21854 4384
rect 21790 4324 21794 4380
rect 21794 4324 21850 4380
rect 21850 4324 21854 4380
rect 21790 4320 21854 4324
rect 21870 4380 21934 4384
rect 21870 4324 21874 4380
rect 21874 4324 21930 4380
rect 21930 4324 21934 4380
rect 21870 4320 21934 4324
rect 21950 4380 22014 4384
rect 21950 4324 21954 4380
rect 21954 4324 22010 4380
rect 22010 4324 22014 4380
rect 21950 4320 22014 4324
rect 22030 4380 22094 4384
rect 22030 4324 22034 4380
rect 22034 4324 22090 4380
rect 22090 4324 22094 4380
rect 22030 4320 22094 4324
rect 28736 4380 28800 4384
rect 28736 4324 28740 4380
rect 28740 4324 28796 4380
rect 28796 4324 28800 4380
rect 28736 4320 28800 4324
rect 28816 4380 28880 4384
rect 28816 4324 28820 4380
rect 28820 4324 28876 4380
rect 28876 4324 28880 4380
rect 28816 4320 28880 4324
rect 28896 4380 28960 4384
rect 28896 4324 28900 4380
rect 28900 4324 28956 4380
rect 28956 4324 28960 4380
rect 28896 4320 28960 4324
rect 28976 4380 29040 4384
rect 28976 4324 28980 4380
rect 28980 4324 29036 4380
rect 29036 4324 29040 4380
rect 28976 4320 29040 4324
rect 4425 3836 4489 3840
rect 4425 3780 4429 3836
rect 4429 3780 4485 3836
rect 4485 3780 4489 3836
rect 4425 3776 4489 3780
rect 4505 3836 4569 3840
rect 4505 3780 4509 3836
rect 4509 3780 4565 3836
rect 4565 3780 4569 3836
rect 4505 3776 4569 3780
rect 4585 3836 4649 3840
rect 4585 3780 4589 3836
rect 4589 3780 4645 3836
rect 4645 3780 4649 3836
rect 4585 3776 4649 3780
rect 4665 3836 4729 3840
rect 4665 3780 4669 3836
rect 4669 3780 4725 3836
rect 4725 3780 4729 3836
rect 4665 3776 4729 3780
rect 11371 3836 11435 3840
rect 11371 3780 11375 3836
rect 11375 3780 11431 3836
rect 11431 3780 11435 3836
rect 11371 3776 11435 3780
rect 11451 3836 11515 3840
rect 11451 3780 11455 3836
rect 11455 3780 11511 3836
rect 11511 3780 11515 3836
rect 11451 3776 11515 3780
rect 11531 3836 11595 3840
rect 11531 3780 11535 3836
rect 11535 3780 11591 3836
rect 11591 3780 11595 3836
rect 11531 3776 11595 3780
rect 11611 3836 11675 3840
rect 11611 3780 11615 3836
rect 11615 3780 11671 3836
rect 11671 3780 11675 3836
rect 11611 3776 11675 3780
rect 18317 3836 18381 3840
rect 18317 3780 18321 3836
rect 18321 3780 18377 3836
rect 18377 3780 18381 3836
rect 18317 3776 18381 3780
rect 18397 3836 18461 3840
rect 18397 3780 18401 3836
rect 18401 3780 18457 3836
rect 18457 3780 18461 3836
rect 18397 3776 18461 3780
rect 18477 3836 18541 3840
rect 18477 3780 18481 3836
rect 18481 3780 18537 3836
rect 18537 3780 18541 3836
rect 18477 3776 18541 3780
rect 18557 3836 18621 3840
rect 18557 3780 18561 3836
rect 18561 3780 18617 3836
rect 18617 3780 18621 3836
rect 18557 3776 18621 3780
rect 25263 3836 25327 3840
rect 25263 3780 25267 3836
rect 25267 3780 25323 3836
rect 25323 3780 25327 3836
rect 25263 3776 25327 3780
rect 25343 3836 25407 3840
rect 25343 3780 25347 3836
rect 25347 3780 25403 3836
rect 25403 3780 25407 3836
rect 25343 3776 25407 3780
rect 25423 3836 25487 3840
rect 25423 3780 25427 3836
rect 25427 3780 25483 3836
rect 25483 3780 25487 3836
rect 25423 3776 25487 3780
rect 25503 3836 25567 3840
rect 25503 3780 25507 3836
rect 25507 3780 25563 3836
rect 25563 3780 25567 3836
rect 25503 3776 25567 3780
rect 7898 3292 7962 3296
rect 7898 3236 7902 3292
rect 7902 3236 7958 3292
rect 7958 3236 7962 3292
rect 7898 3232 7962 3236
rect 7978 3292 8042 3296
rect 7978 3236 7982 3292
rect 7982 3236 8038 3292
rect 8038 3236 8042 3292
rect 7978 3232 8042 3236
rect 8058 3292 8122 3296
rect 8058 3236 8062 3292
rect 8062 3236 8118 3292
rect 8118 3236 8122 3292
rect 8058 3232 8122 3236
rect 8138 3292 8202 3296
rect 8138 3236 8142 3292
rect 8142 3236 8198 3292
rect 8198 3236 8202 3292
rect 8138 3232 8202 3236
rect 14844 3292 14908 3296
rect 14844 3236 14848 3292
rect 14848 3236 14904 3292
rect 14904 3236 14908 3292
rect 14844 3232 14908 3236
rect 14924 3292 14988 3296
rect 14924 3236 14928 3292
rect 14928 3236 14984 3292
rect 14984 3236 14988 3292
rect 14924 3232 14988 3236
rect 15004 3292 15068 3296
rect 15004 3236 15008 3292
rect 15008 3236 15064 3292
rect 15064 3236 15068 3292
rect 15004 3232 15068 3236
rect 15084 3292 15148 3296
rect 15084 3236 15088 3292
rect 15088 3236 15144 3292
rect 15144 3236 15148 3292
rect 15084 3232 15148 3236
rect 21790 3292 21854 3296
rect 21790 3236 21794 3292
rect 21794 3236 21850 3292
rect 21850 3236 21854 3292
rect 21790 3232 21854 3236
rect 21870 3292 21934 3296
rect 21870 3236 21874 3292
rect 21874 3236 21930 3292
rect 21930 3236 21934 3292
rect 21870 3232 21934 3236
rect 21950 3292 22014 3296
rect 21950 3236 21954 3292
rect 21954 3236 22010 3292
rect 22010 3236 22014 3292
rect 21950 3232 22014 3236
rect 22030 3292 22094 3296
rect 22030 3236 22034 3292
rect 22034 3236 22090 3292
rect 22090 3236 22094 3292
rect 22030 3232 22094 3236
rect 28736 3292 28800 3296
rect 28736 3236 28740 3292
rect 28740 3236 28796 3292
rect 28796 3236 28800 3292
rect 28736 3232 28800 3236
rect 28816 3292 28880 3296
rect 28816 3236 28820 3292
rect 28820 3236 28876 3292
rect 28876 3236 28880 3292
rect 28816 3232 28880 3236
rect 28896 3292 28960 3296
rect 28896 3236 28900 3292
rect 28900 3236 28956 3292
rect 28956 3236 28960 3292
rect 28896 3232 28960 3236
rect 28976 3292 29040 3296
rect 28976 3236 28980 3292
rect 28980 3236 29036 3292
rect 29036 3236 29040 3292
rect 28976 3232 29040 3236
rect 4425 2748 4489 2752
rect 4425 2692 4429 2748
rect 4429 2692 4485 2748
rect 4485 2692 4489 2748
rect 4425 2688 4489 2692
rect 4505 2748 4569 2752
rect 4505 2692 4509 2748
rect 4509 2692 4565 2748
rect 4565 2692 4569 2748
rect 4505 2688 4569 2692
rect 4585 2748 4649 2752
rect 4585 2692 4589 2748
rect 4589 2692 4645 2748
rect 4645 2692 4649 2748
rect 4585 2688 4649 2692
rect 4665 2748 4729 2752
rect 4665 2692 4669 2748
rect 4669 2692 4725 2748
rect 4725 2692 4729 2748
rect 4665 2688 4729 2692
rect 11371 2748 11435 2752
rect 11371 2692 11375 2748
rect 11375 2692 11431 2748
rect 11431 2692 11435 2748
rect 11371 2688 11435 2692
rect 11451 2748 11515 2752
rect 11451 2692 11455 2748
rect 11455 2692 11511 2748
rect 11511 2692 11515 2748
rect 11451 2688 11515 2692
rect 11531 2748 11595 2752
rect 11531 2692 11535 2748
rect 11535 2692 11591 2748
rect 11591 2692 11595 2748
rect 11531 2688 11595 2692
rect 11611 2748 11675 2752
rect 11611 2692 11615 2748
rect 11615 2692 11671 2748
rect 11671 2692 11675 2748
rect 11611 2688 11675 2692
rect 18317 2748 18381 2752
rect 18317 2692 18321 2748
rect 18321 2692 18377 2748
rect 18377 2692 18381 2748
rect 18317 2688 18381 2692
rect 18397 2748 18461 2752
rect 18397 2692 18401 2748
rect 18401 2692 18457 2748
rect 18457 2692 18461 2748
rect 18397 2688 18461 2692
rect 18477 2748 18541 2752
rect 18477 2692 18481 2748
rect 18481 2692 18537 2748
rect 18537 2692 18541 2748
rect 18477 2688 18541 2692
rect 18557 2748 18621 2752
rect 18557 2692 18561 2748
rect 18561 2692 18617 2748
rect 18617 2692 18621 2748
rect 18557 2688 18621 2692
rect 25263 2748 25327 2752
rect 25263 2692 25267 2748
rect 25267 2692 25323 2748
rect 25323 2692 25327 2748
rect 25263 2688 25327 2692
rect 25343 2748 25407 2752
rect 25343 2692 25347 2748
rect 25347 2692 25403 2748
rect 25403 2692 25407 2748
rect 25343 2688 25407 2692
rect 25423 2748 25487 2752
rect 25423 2692 25427 2748
rect 25427 2692 25483 2748
rect 25483 2692 25487 2748
rect 25423 2688 25487 2692
rect 25503 2748 25567 2752
rect 25503 2692 25507 2748
rect 25507 2692 25563 2748
rect 25563 2692 25567 2748
rect 25503 2688 25567 2692
rect 7898 2204 7962 2208
rect 7898 2148 7902 2204
rect 7902 2148 7958 2204
rect 7958 2148 7962 2204
rect 7898 2144 7962 2148
rect 7978 2204 8042 2208
rect 7978 2148 7982 2204
rect 7982 2148 8038 2204
rect 8038 2148 8042 2204
rect 7978 2144 8042 2148
rect 8058 2204 8122 2208
rect 8058 2148 8062 2204
rect 8062 2148 8118 2204
rect 8118 2148 8122 2204
rect 8058 2144 8122 2148
rect 8138 2204 8202 2208
rect 8138 2148 8142 2204
rect 8142 2148 8198 2204
rect 8198 2148 8202 2204
rect 8138 2144 8202 2148
rect 14844 2204 14908 2208
rect 14844 2148 14848 2204
rect 14848 2148 14904 2204
rect 14904 2148 14908 2204
rect 14844 2144 14908 2148
rect 14924 2204 14988 2208
rect 14924 2148 14928 2204
rect 14928 2148 14984 2204
rect 14984 2148 14988 2204
rect 14924 2144 14988 2148
rect 15004 2204 15068 2208
rect 15004 2148 15008 2204
rect 15008 2148 15064 2204
rect 15064 2148 15068 2204
rect 15004 2144 15068 2148
rect 15084 2204 15148 2208
rect 15084 2148 15088 2204
rect 15088 2148 15144 2204
rect 15144 2148 15148 2204
rect 15084 2144 15148 2148
rect 21790 2204 21854 2208
rect 21790 2148 21794 2204
rect 21794 2148 21850 2204
rect 21850 2148 21854 2204
rect 21790 2144 21854 2148
rect 21870 2204 21934 2208
rect 21870 2148 21874 2204
rect 21874 2148 21930 2204
rect 21930 2148 21934 2204
rect 21870 2144 21934 2148
rect 21950 2204 22014 2208
rect 21950 2148 21954 2204
rect 21954 2148 22010 2204
rect 22010 2148 22014 2204
rect 21950 2144 22014 2148
rect 22030 2204 22094 2208
rect 22030 2148 22034 2204
rect 22034 2148 22090 2204
rect 22090 2148 22094 2204
rect 22030 2144 22094 2148
rect 28736 2204 28800 2208
rect 28736 2148 28740 2204
rect 28740 2148 28796 2204
rect 28796 2148 28800 2204
rect 28736 2144 28800 2148
rect 28816 2204 28880 2208
rect 28816 2148 28820 2204
rect 28820 2148 28876 2204
rect 28876 2148 28880 2204
rect 28816 2144 28880 2148
rect 28896 2204 28960 2208
rect 28896 2148 28900 2204
rect 28900 2148 28956 2204
rect 28956 2148 28960 2204
rect 28896 2144 28960 2148
rect 28976 2204 29040 2208
rect 28976 2148 28980 2204
rect 28980 2148 29036 2204
rect 29036 2148 29040 2204
rect 28976 2144 29040 2148
rect 12756 1396 12820 1460
<< metal4 >>
rect 16435 31788 16501 31789
rect 16435 31724 16436 31788
rect 16500 31724 16501 31788
rect 16435 31723 16501 31724
rect 4417 31040 4737 31600
rect 4417 30976 4425 31040
rect 4489 30976 4505 31040
rect 4569 30976 4585 31040
rect 4649 30976 4665 31040
rect 4729 30976 4737 31040
rect 4417 29952 4737 30976
rect 7890 31584 8210 31600
rect 7890 31520 7898 31584
rect 7962 31520 7978 31584
rect 8042 31520 8058 31584
rect 8122 31520 8138 31584
rect 8202 31520 8210 31584
rect 7890 30496 8210 31520
rect 7890 30432 7898 30496
rect 7962 30432 7978 30496
rect 8042 30432 8058 30496
rect 8122 30432 8138 30496
rect 8202 30432 8210 30496
rect 6867 30428 6933 30429
rect 6867 30364 6868 30428
rect 6932 30364 6933 30428
rect 6867 30363 6933 30364
rect 4417 29888 4425 29952
rect 4489 29888 4505 29952
rect 4569 29888 4585 29952
rect 4649 29888 4665 29952
rect 4729 29888 4737 29952
rect 4417 28864 4737 29888
rect 4417 28800 4425 28864
rect 4489 28800 4505 28864
rect 4569 28800 4585 28864
rect 4649 28800 4665 28864
rect 4729 28800 4737 28864
rect 4417 27776 4737 28800
rect 4417 27712 4425 27776
rect 4489 27712 4505 27776
rect 4569 27712 4585 27776
rect 4649 27712 4665 27776
rect 4729 27712 4737 27776
rect 4417 26688 4737 27712
rect 6870 27437 6930 30363
rect 7890 29408 8210 30432
rect 7890 29344 7898 29408
rect 7962 29344 7978 29408
rect 8042 29344 8058 29408
rect 8122 29344 8138 29408
rect 8202 29344 8210 29408
rect 7890 28320 8210 29344
rect 7890 28256 7898 28320
rect 7962 28256 7978 28320
rect 8042 28256 8058 28320
rect 8122 28256 8138 28320
rect 8202 28256 8210 28320
rect 6867 27436 6933 27437
rect 6867 27372 6868 27436
rect 6932 27372 6933 27436
rect 6867 27371 6933 27372
rect 4417 26624 4425 26688
rect 4489 26624 4505 26688
rect 4569 26624 4585 26688
rect 4649 26624 4665 26688
rect 4729 26624 4737 26688
rect 4417 25600 4737 26624
rect 4417 25536 4425 25600
rect 4489 25536 4505 25600
rect 4569 25536 4585 25600
rect 4649 25536 4665 25600
rect 4729 25536 4737 25600
rect 4417 24512 4737 25536
rect 4417 24448 4425 24512
rect 4489 24448 4505 24512
rect 4569 24448 4585 24512
rect 4649 24448 4665 24512
rect 4729 24448 4737 24512
rect 4417 23424 4737 24448
rect 4417 23360 4425 23424
rect 4489 23360 4505 23424
rect 4569 23360 4585 23424
rect 4649 23360 4665 23424
rect 4729 23360 4737 23424
rect 4417 22336 4737 23360
rect 4417 22272 4425 22336
rect 4489 22272 4505 22336
rect 4569 22272 4585 22336
rect 4649 22272 4665 22336
rect 4729 22272 4737 22336
rect 4417 21248 4737 22272
rect 4417 21184 4425 21248
rect 4489 21184 4505 21248
rect 4569 21184 4585 21248
rect 4649 21184 4665 21248
rect 4729 21184 4737 21248
rect 4417 20160 4737 21184
rect 4417 20096 4425 20160
rect 4489 20096 4505 20160
rect 4569 20096 4585 20160
rect 4649 20096 4665 20160
rect 4729 20096 4737 20160
rect 4417 19072 4737 20096
rect 4417 19008 4425 19072
rect 4489 19008 4505 19072
rect 4569 19008 4585 19072
rect 4649 19008 4665 19072
rect 4729 19008 4737 19072
rect 4417 17984 4737 19008
rect 4417 17920 4425 17984
rect 4489 17920 4505 17984
rect 4569 17920 4585 17984
rect 4649 17920 4665 17984
rect 4729 17920 4737 17984
rect 4417 16896 4737 17920
rect 4417 16832 4425 16896
rect 4489 16832 4505 16896
rect 4569 16832 4585 16896
rect 4649 16832 4665 16896
rect 4729 16832 4737 16896
rect 4417 15808 4737 16832
rect 4417 15744 4425 15808
rect 4489 15744 4505 15808
rect 4569 15744 4585 15808
rect 4649 15744 4665 15808
rect 4729 15744 4737 15808
rect 4417 14720 4737 15744
rect 4417 14656 4425 14720
rect 4489 14656 4505 14720
rect 4569 14656 4585 14720
rect 4649 14656 4665 14720
rect 4729 14656 4737 14720
rect 4417 13632 4737 14656
rect 4417 13568 4425 13632
rect 4489 13568 4505 13632
rect 4569 13568 4585 13632
rect 4649 13568 4665 13632
rect 4729 13568 4737 13632
rect 4417 12544 4737 13568
rect 4417 12480 4425 12544
rect 4489 12480 4505 12544
rect 4569 12480 4585 12544
rect 4649 12480 4665 12544
rect 4729 12480 4737 12544
rect 4417 11456 4737 12480
rect 4417 11392 4425 11456
rect 4489 11392 4505 11456
rect 4569 11392 4585 11456
rect 4649 11392 4665 11456
rect 4729 11392 4737 11456
rect 4417 10368 4737 11392
rect 4417 10304 4425 10368
rect 4489 10304 4505 10368
rect 4569 10304 4585 10368
rect 4649 10304 4665 10368
rect 4729 10304 4737 10368
rect 4417 9280 4737 10304
rect 4417 9216 4425 9280
rect 4489 9216 4505 9280
rect 4569 9216 4585 9280
rect 4649 9216 4665 9280
rect 4729 9216 4737 9280
rect 4417 8192 4737 9216
rect 4417 8128 4425 8192
rect 4489 8128 4505 8192
rect 4569 8128 4585 8192
rect 4649 8128 4665 8192
rect 4729 8128 4737 8192
rect 4417 7104 4737 8128
rect 4417 7040 4425 7104
rect 4489 7040 4505 7104
rect 4569 7040 4585 7104
rect 4649 7040 4665 7104
rect 4729 7040 4737 7104
rect 4417 6016 4737 7040
rect 4417 5952 4425 6016
rect 4489 5952 4505 6016
rect 4569 5952 4585 6016
rect 4649 5952 4665 6016
rect 4729 5952 4737 6016
rect 4417 4928 4737 5952
rect 4417 4864 4425 4928
rect 4489 4864 4505 4928
rect 4569 4864 4585 4928
rect 4649 4864 4665 4928
rect 4729 4864 4737 4928
rect 4417 3840 4737 4864
rect 4417 3776 4425 3840
rect 4489 3776 4505 3840
rect 4569 3776 4585 3840
rect 4649 3776 4665 3840
rect 4729 3776 4737 3840
rect 4417 2752 4737 3776
rect 4417 2688 4425 2752
rect 4489 2688 4505 2752
rect 4569 2688 4585 2752
rect 4649 2688 4665 2752
rect 4729 2688 4737 2752
rect 4417 2128 4737 2688
rect 7890 27232 8210 28256
rect 7890 27168 7898 27232
rect 7962 27168 7978 27232
rect 8042 27168 8058 27232
rect 8122 27168 8138 27232
rect 8202 27168 8210 27232
rect 7890 26144 8210 27168
rect 7890 26080 7898 26144
rect 7962 26080 7978 26144
rect 8042 26080 8058 26144
rect 8122 26080 8138 26144
rect 8202 26080 8210 26144
rect 7890 25056 8210 26080
rect 7890 24992 7898 25056
rect 7962 24992 7978 25056
rect 8042 24992 8058 25056
rect 8122 24992 8138 25056
rect 8202 24992 8210 25056
rect 7890 23968 8210 24992
rect 7890 23904 7898 23968
rect 7962 23904 7978 23968
rect 8042 23904 8058 23968
rect 8122 23904 8138 23968
rect 8202 23904 8210 23968
rect 7890 22880 8210 23904
rect 7890 22816 7898 22880
rect 7962 22816 7978 22880
rect 8042 22816 8058 22880
rect 8122 22816 8138 22880
rect 8202 22816 8210 22880
rect 7890 21792 8210 22816
rect 7890 21728 7898 21792
rect 7962 21728 7978 21792
rect 8042 21728 8058 21792
rect 8122 21728 8138 21792
rect 8202 21728 8210 21792
rect 7890 20704 8210 21728
rect 7890 20640 7898 20704
rect 7962 20640 7978 20704
rect 8042 20640 8058 20704
rect 8122 20640 8138 20704
rect 8202 20640 8210 20704
rect 7890 19616 8210 20640
rect 7890 19552 7898 19616
rect 7962 19552 7978 19616
rect 8042 19552 8058 19616
rect 8122 19552 8138 19616
rect 8202 19552 8210 19616
rect 7890 18528 8210 19552
rect 7890 18464 7898 18528
rect 7962 18464 7978 18528
rect 8042 18464 8058 18528
rect 8122 18464 8138 18528
rect 8202 18464 8210 18528
rect 7890 17440 8210 18464
rect 7890 17376 7898 17440
rect 7962 17376 7978 17440
rect 8042 17376 8058 17440
rect 8122 17376 8138 17440
rect 8202 17376 8210 17440
rect 7890 16352 8210 17376
rect 7890 16288 7898 16352
rect 7962 16288 7978 16352
rect 8042 16288 8058 16352
rect 8122 16288 8138 16352
rect 8202 16288 8210 16352
rect 7890 15264 8210 16288
rect 7890 15200 7898 15264
rect 7962 15200 7978 15264
rect 8042 15200 8058 15264
rect 8122 15200 8138 15264
rect 8202 15200 8210 15264
rect 7890 14176 8210 15200
rect 7890 14112 7898 14176
rect 7962 14112 7978 14176
rect 8042 14112 8058 14176
rect 8122 14112 8138 14176
rect 8202 14112 8210 14176
rect 7890 13088 8210 14112
rect 7890 13024 7898 13088
rect 7962 13024 7978 13088
rect 8042 13024 8058 13088
rect 8122 13024 8138 13088
rect 8202 13024 8210 13088
rect 7890 12000 8210 13024
rect 7890 11936 7898 12000
rect 7962 11936 7978 12000
rect 8042 11936 8058 12000
rect 8122 11936 8138 12000
rect 8202 11936 8210 12000
rect 7890 10912 8210 11936
rect 7890 10848 7898 10912
rect 7962 10848 7978 10912
rect 8042 10848 8058 10912
rect 8122 10848 8138 10912
rect 8202 10848 8210 10912
rect 7890 9824 8210 10848
rect 7890 9760 7898 9824
rect 7962 9760 7978 9824
rect 8042 9760 8058 9824
rect 8122 9760 8138 9824
rect 8202 9760 8210 9824
rect 7890 8736 8210 9760
rect 7890 8672 7898 8736
rect 7962 8672 7978 8736
rect 8042 8672 8058 8736
rect 8122 8672 8138 8736
rect 8202 8672 8210 8736
rect 7890 7648 8210 8672
rect 7890 7584 7898 7648
rect 7962 7584 7978 7648
rect 8042 7584 8058 7648
rect 8122 7584 8138 7648
rect 8202 7584 8210 7648
rect 7890 6560 8210 7584
rect 7890 6496 7898 6560
rect 7962 6496 7978 6560
rect 8042 6496 8058 6560
rect 8122 6496 8138 6560
rect 8202 6496 8210 6560
rect 7890 5472 8210 6496
rect 7890 5408 7898 5472
rect 7962 5408 7978 5472
rect 8042 5408 8058 5472
rect 8122 5408 8138 5472
rect 8202 5408 8210 5472
rect 7890 4384 8210 5408
rect 7890 4320 7898 4384
rect 7962 4320 7978 4384
rect 8042 4320 8058 4384
rect 8122 4320 8138 4384
rect 8202 4320 8210 4384
rect 7890 3296 8210 4320
rect 7890 3232 7898 3296
rect 7962 3232 7978 3296
rect 8042 3232 8058 3296
rect 8122 3232 8138 3296
rect 8202 3232 8210 3296
rect 7890 2208 8210 3232
rect 7890 2144 7898 2208
rect 7962 2144 7978 2208
rect 8042 2144 8058 2208
rect 8122 2144 8138 2208
rect 8202 2144 8210 2208
rect 7890 2128 8210 2144
rect 11363 31040 11683 31600
rect 11363 30976 11371 31040
rect 11435 30976 11451 31040
rect 11515 30976 11531 31040
rect 11595 30976 11611 31040
rect 11675 30976 11683 31040
rect 11363 29952 11683 30976
rect 14836 31584 15156 31600
rect 14836 31520 14844 31584
rect 14908 31520 14924 31584
rect 14988 31520 15004 31584
rect 15068 31520 15084 31584
rect 15148 31520 15156 31584
rect 14836 30496 15156 31520
rect 15331 31380 15397 31381
rect 15331 31316 15332 31380
rect 15396 31316 15397 31380
rect 15331 31315 15397 31316
rect 14836 30432 14844 30496
rect 14908 30432 14924 30496
rect 14988 30432 15004 30496
rect 15068 30432 15084 30496
rect 15148 30432 15156 30496
rect 14595 30156 14661 30157
rect 14595 30092 14596 30156
rect 14660 30092 14661 30156
rect 14595 30091 14661 30092
rect 11363 29888 11371 29952
rect 11435 29888 11451 29952
rect 11515 29888 11531 29952
rect 11595 29888 11611 29952
rect 11675 29888 11683 29952
rect 11363 28864 11683 29888
rect 12939 29612 13005 29613
rect 12939 29548 12940 29612
rect 13004 29548 13005 29612
rect 12939 29547 13005 29548
rect 11363 28800 11371 28864
rect 11435 28800 11451 28864
rect 11515 28800 11531 28864
rect 11595 28800 11611 28864
rect 11675 28800 11683 28864
rect 11363 27776 11683 28800
rect 12755 27980 12821 27981
rect 12755 27916 12756 27980
rect 12820 27916 12821 27980
rect 12755 27915 12821 27916
rect 11363 27712 11371 27776
rect 11435 27712 11451 27776
rect 11515 27712 11531 27776
rect 11595 27712 11611 27776
rect 11675 27712 11683 27776
rect 11363 26688 11683 27712
rect 11363 26624 11371 26688
rect 11435 26624 11451 26688
rect 11515 26624 11531 26688
rect 11595 26624 11611 26688
rect 11675 26624 11683 26688
rect 11363 25600 11683 26624
rect 11363 25536 11371 25600
rect 11435 25536 11451 25600
rect 11515 25536 11531 25600
rect 11595 25536 11611 25600
rect 11675 25536 11683 25600
rect 11363 24512 11683 25536
rect 11363 24448 11371 24512
rect 11435 24448 11451 24512
rect 11515 24448 11531 24512
rect 11595 24448 11611 24512
rect 11675 24448 11683 24512
rect 11363 23424 11683 24448
rect 11363 23360 11371 23424
rect 11435 23360 11451 23424
rect 11515 23360 11531 23424
rect 11595 23360 11611 23424
rect 11675 23360 11683 23424
rect 11363 22336 11683 23360
rect 11363 22272 11371 22336
rect 11435 22272 11451 22336
rect 11515 22272 11531 22336
rect 11595 22272 11611 22336
rect 11675 22272 11683 22336
rect 11363 21248 11683 22272
rect 11363 21184 11371 21248
rect 11435 21184 11451 21248
rect 11515 21184 11531 21248
rect 11595 21184 11611 21248
rect 11675 21184 11683 21248
rect 11363 20160 11683 21184
rect 11363 20096 11371 20160
rect 11435 20096 11451 20160
rect 11515 20096 11531 20160
rect 11595 20096 11611 20160
rect 11675 20096 11683 20160
rect 11363 19072 11683 20096
rect 11363 19008 11371 19072
rect 11435 19008 11451 19072
rect 11515 19008 11531 19072
rect 11595 19008 11611 19072
rect 11675 19008 11683 19072
rect 11363 17984 11683 19008
rect 11363 17920 11371 17984
rect 11435 17920 11451 17984
rect 11515 17920 11531 17984
rect 11595 17920 11611 17984
rect 11675 17920 11683 17984
rect 11363 16896 11683 17920
rect 11363 16832 11371 16896
rect 11435 16832 11451 16896
rect 11515 16832 11531 16896
rect 11595 16832 11611 16896
rect 11675 16832 11683 16896
rect 11363 15808 11683 16832
rect 11363 15744 11371 15808
rect 11435 15744 11451 15808
rect 11515 15744 11531 15808
rect 11595 15744 11611 15808
rect 11675 15744 11683 15808
rect 11363 14720 11683 15744
rect 11363 14656 11371 14720
rect 11435 14656 11451 14720
rect 11515 14656 11531 14720
rect 11595 14656 11611 14720
rect 11675 14656 11683 14720
rect 11363 13632 11683 14656
rect 11363 13568 11371 13632
rect 11435 13568 11451 13632
rect 11515 13568 11531 13632
rect 11595 13568 11611 13632
rect 11675 13568 11683 13632
rect 11363 12544 11683 13568
rect 11363 12480 11371 12544
rect 11435 12480 11451 12544
rect 11515 12480 11531 12544
rect 11595 12480 11611 12544
rect 11675 12480 11683 12544
rect 11363 11456 11683 12480
rect 11363 11392 11371 11456
rect 11435 11392 11451 11456
rect 11515 11392 11531 11456
rect 11595 11392 11611 11456
rect 11675 11392 11683 11456
rect 11363 10368 11683 11392
rect 11363 10304 11371 10368
rect 11435 10304 11451 10368
rect 11515 10304 11531 10368
rect 11595 10304 11611 10368
rect 11675 10304 11683 10368
rect 11363 9280 11683 10304
rect 11363 9216 11371 9280
rect 11435 9216 11451 9280
rect 11515 9216 11531 9280
rect 11595 9216 11611 9280
rect 11675 9216 11683 9280
rect 11363 8192 11683 9216
rect 11363 8128 11371 8192
rect 11435 8128 11451 8192
rect 11515 8128 11531 8192
rect 11595 8128 11611 8192
rect 11675 8128 11683 8192
rect 11363 7104 11683 8128
rect 11363 7040 11371 7104
rect 11435 7040 11451 7104
rect 11515 7040 11531 7104
rect 11595 7040 11611 7104
rect 11675 7040 11683 7104
rect 11363 6016 11683 7040
rect 11363 5952 11371 6016
rect 11435 5952 11451 6016
rect 11515 5952 11531 6016
rect 11595 5952 11611 6016
rect 11675 5952 11683 6016
rect 11363 4928 11683 5952
rect 11363 4864 11371 4928
rect 11435 4864 11451 4928
rect 11515 4864 11531 4928
rect 11595 4864 11611 4928
rect 11675 4864 11683 4928
rect 11363 3840 11683 4864
rect 11363 3776 11371 3840
rect 11435 3776 11451 3840
rect 11515 3776 11531 3840
rect 11595 3776 11611 3840
rect 11675 3776 11683 3840
rect 11363 2752 11683 3776
rect 11363 2688 11371 2752
rect 11435 2688 11451 2752
rect 11515 2688 11531 2752
rect 11595 2688 11611 2752
rect 11675 2688 11683 2752
rect 11363 2128 11683 2688
rect 12758 1461 12818 27915
rect 12942 27301 13002 29547
rect 12939 27300 13005 27301
rect 12939 27236 12940 27300
rect 13004 27236 13005 27300
rect 12939 27235 13005 27236
rect 14598 26485 14658 30091
rect 14836 29408 15156 30432
rect 15334 29749 15394 31315
rect 15331 29748 15397 29749
rect 15331 29684 15332 29748
rect 15396 29684 15397 29748
rect 15331 29683 15397 29684
rect 15699 29748 15765 29749
rect 15699 29684 15700 29748
rect 15764 29684 15765 29748
rect 15699 29683 15765 29684
rect 14836 29344 14844 29408
rect 14908 29344 14924 29408
rect 14988 29344 15004 29408
rect 15068 29344 15084 29408
rect 15148 29344 15156 29408
rect 14836 28320 15156 29344
rect 15702 29205 15762 29683
rect 16438 29205 16498 31723
rect 18309 31040 18629 31600
rect 18309 30976 18317 31040
rect 18381 30976 18397 31040
rect 18461 30976 18477 31040
rect 18541 30976 18557 31040
rect 18621 30976 18629 31040
rect 16619 30428 16685 30429
rect 16619 30364 16620 30428
rect 16684 30364 16685 30428
rect 16619 30363 16685 30364
rect 16622 29477 16682 30363
rect 18309 29952 18629 30976
rect 18309 29888 18317 29952
rect 18381 29888 18397 29952
rect 18461 29888 18477 29952
rect 18541 29888 18557 29952
rect 18621 29888 18629 29952
rect 16619 29476 16685 29477
rect 16619 29412 16620 29476
rect 16684 29412 16685 29476
rect 16619 29411 16685 29412
rect 15699 29204 15765 29205
rect 15699 29140 15700 29204
rect 15764 29140 15765 29204
rect 15699 29139 15765 29140
rect 16435 29204 16501 29205
rect 16435 29140 16436 29204
rect 16500 29140 16501 29204
rect 16435 29139 16501 29140
rect 14836 28256 14844 28320
rect 14908 28256 14924 28320
rect 14988 28256 15004 28320
rect 15068 28256 15084 28320
rect 15148 28256 15156 28320
rect 14836 27232 15156 28256
rect 14836 27168 14844 27232
rect 14908 27168 14924 27232
rect 14988 27168 15004 27232
rect 15068 27168 15084 27232
rect 15148 27168 15156 27232
rect 14595 26484 14661 26485
rect 14595 26420 14596 26484
rect 14660 26420 14661 26484
rect 14595 26419 14661 26420
rect 14836 26144 15156 27168
rect 14836 26080 14844 26144
rect 14908 26080 14924 26144
rect 14988 26080 15004 26144
rect 15068 26080 15084 26144
rect 15148 26080 15156 26144
rect 14836 25056 15156 26080
rect 14836 24992 14844 25056
rect 14908 24992 14924 25056
rect 14988 24992 15004 25056
rect 15068 24992 15084 25056
rect 15148 24992 15156 25056
rect 14836 23968 15156 24992
rect 14836 23904 14844 23968
rect 14908 23904 14924 23968
rect 14988 23904 15004 23968
rect 15068 23904 15084 23968
rect 15148 23904 15156 23968
rect 14836 22880 15156 23904
rect 14836 22816 14844 22880
rect 14908 22816 14924 22880
rect 14988 22816 15004 22880
rect 15068 22816 15084 22880
rect 15148 22816 15156 22880
rect 14836 21792 15156 22816
rect 14836 21728 14844 21792
rect 14908 21728 14924 21792
rect 14988 21728 15004 21792
rect 15068 21728 15084 21792
rect 15148 21728 15156 21792
rect 14836 20704 15156 21728
rect 14836 20640 14844 20704
rect 14908 20640 14924 20704
rect 14988 20640 15004 20704
rect 15068 20640 15084 20704
rect 15148 20640 15156 20704
rect 14836 19616 15156 20640
rect 14836 19552 14844 19616
rect 14908 19552 14924 19616
rect 14988 19552 15004 19616
rect 15068 19552 15084 19616
rect 15148 19552 15156 19616
rect 14836 18528 15156 19552
rect 14836 18464 14844 18528
rect 14908 18464 14924 18528
rect 14988 18464 15004 18528
rect 15068 18464 15084 18528
rect 15148 18464 15156 18528
rect 14836 17440 15156 18464
rect 14836 17376 14844 17440
rect 14908 17376 14924 17440
rect 14988 17376 15004 17440
rect 15068 17376 15084 17440
rect 15148 17376 15156 17440
rect 14836 16352 15156 17376
rect 14836 16288 14844 16352
rect 14908 16288 14924 16352
rect 14988 16288 15004 16352
rect 15068 16288 15084 16352
rect 15148 16288 15156 16352
rect 14836 15264 15156 16288
rect 14836 15200 14844 15264
rect 14908 15200 14924 15264
rect 14988 15200 15004 15264
rect 15068 15200 15084 15264
rect 15148 15200 15156 15264
rect 14836 14176 15156 15200
rect 14836 14112 14844 14176
rect 14908 14112 14924 14176
rect 14988 14112 15004 14176
rect 15068 14112 15084 14176
rect 15148 14112 15156 14176
rect 14836 13088 15156 14112
rect 14836 13024 14844 13088
rect 14908 13024 14924 13088
rect 14988 13024 15004 13088
rect 15068 13024 15084 13088
rect 15148 13024 15156 13088
rect 14836 12000 15156 13024
rect 14836 11936 14844 12000
rect 14908 11936 14924 12000
rect 14988 11936 15004 12000
rect 15068 11936 15084 12000
rect 15148 11936 15156 12000
rect 14836 10912 15156 11936
rect 14836 10848 14844 10912
rect 14908 10848 14924 10912
rect 14988 10848 15004 10912
rect 15068 10848 15084 10912
rect 15148 10848 15156 10912
rect 14836 9824 15156 10848
rect 14836 9760 14844 9824
rect 14908 9760 14924 9824
rect 14988 9760 15004 9824
rect 15068 9760 15084 9824
rect 15148 9760 15156 9824
rect 14836 8736 15156 9760
rect 14836 8672 14844 8736
rect 14908 8672 14924 8736
rect 14988 8672 15004 8736
rect 15068 8672 15084 8736
rect 15148 8672 15156 8736
rect 14836 7648 15156 8672
rect 14836 7584 14844 7648
rect 14908 7584 14924 7648
rect 14988 7584 15004 7648
rect 15068 7584 15084 7648
rect 15148 7584 15156 7648
rect 14836 6560 15156 7584
rect 14836 6496 14844 6560
rect 14908 6496 14924 6560
rect 14988 6496 15004 6560
rect 15068 6496 15084 6560
rect 15148 6496 15156 6560
rect 14836 5472 15156 6496
rect 14836 5408 14844 5472
rect 14908 5408 14924 5472
rect 14988 5408 15004 5472
rect 15068 5408 15084 5472
rect 15148 5408 15156 5472
rect 14836 4384 15156 5408
rect 14836 4320 14844 4384
rect 14908 4320 14924 4384
rect 14988 4320 15004 4384
rect 15068 4320 15084 4384
rect 15148 4320 15156 4384
rect 14836 3296 15156 4320
rect 14836 3232 14844 3296
rect 14908 3232 14924 3296
rect 14988 3232 15004 3296
rect 15068 3232 15084 3296
rect 15148 3232 15156 3296
rect 14836 2208 15156 3232
rect 14836 2144 14844 2208
rect 14908 2144 14924 2208
rect 14988 2144 15004 2208
rect 15068 2144 15084 2208
rect 15148 2144 15156 2208
rect 14836 2128 15156 2144
rect 18309 28864 18629 29888
rect 18309 28800 18317 28864
rect 18381 28800 18397 28864
rect 18461 28800 18477 28864
rect 18541 28800 18557 28864
rect 18621 28800 18629 28864
rect 18309 27776 18629 28800
rect 18309 27712 18317 27776
rect 18381 27712 18397 27776
rect 18461 27712 18477 27776
rect 18541 27712 18557 27776
rect 18621 27712 18629 27776
rect 18309 26688 18629 27712
rect 18309 26624 18317 26688
rect 18381 26624 18397 26688
rect 18461 26624 18477 26688
rect 18541 26624 18557 26688
rect 18621 26624 18629 26688
rect 18309 25600 18629 26624
rect 18309 25536 18317 25600
rect 18381 25536 18397 25600
rect 18461 25536 18477 25600
rect 18541 25536 18557 25600
rect 18621 25536 18629 25600
rect 18309 24512 18629 25536
rect 18309 24448 18317 24512
rect 18381 24448 18397 24512
rect 18461 24448 18477 24512
rect 18541 24448 18557 24512
rect 18621 24448 18629 24512
rect 18309 23424 18629 24448
rect 18309 23360 18317 23424
rect 18381 23360 18397 23424
rect 18461 23360 18477 23424
rect 18541 23360 18557 23424
rect 18621 23360 18629 23424
rect 18309 22336 18629 23360
rect 18309 22272 18317 22336
rect 18381 22272 18397 22336
rect 18461 22272 18477 22336
rect 18541 22272 18557 22336
rect 18621 22272 18629 22336
rect 18309 21248 18629 22272
rect 18309 21184 18317 21248
rect 18381 21184 18397 21248
rect 18461 21184 18477 21248
rect 18541 21184 18557 21248
rect 18621 21184 18629 21248
rect 18309 20160 18629 21184
rect 18309 20096 18317 20160
rect 18381 20096 18397 20160
rect 18461 20096 18477 20160
rect 18541 20096 18557 20160
rect 18621 20096 18629 20160
rect 18309 19072 18629 20096
rect 18309 19008 18317 19072
rect 18381 19008 18397 19072
rect 18461 19008 18477 19072
rect 18541 19008 18557 19072
rect 18621 19008 18629 19072
rect 18309 17984 18629 19008
rect 18309 17920 18317 17984
rect 18381 17920 18397 17984
rect 18461 17920 18477 17984
rect 18541 17920 18557 17984
rect 18621 17920 18629 17984
rect 18309 16896 18629 17920
rect 18309 16832 18317 16896
rect 18381 16832 18397 16896
rect 18461 16832 18477 16896
rect 18541 16832 18557 16896
rect 18621 16832 18629 16896
rect 18309 15808 18629 16832
rect 18309 15744 18317 15808
rect 18381 15744 18397 15808
rect 18461 15744 18477 15808
rect 18541 15744 18557 15808
rect 18621 15744 18629 15808
rect 18309 14720 18629 15744
rect 18309 14656 18317 14720
rect 18381 14656 18397 14720
rect 18461 14656 18477 14720
rect 18541 14656 18557 14720
rect 18621 14656 18629 14720
rect 18309 13632 18629 14656
rect 18309 13568 18317 13632
rect 18381 13568 18397 13632
rect 18461 13568 18477 13632
rect 18541 13568 18557 13632
rect 18621 13568 18629 13632
rect 18309 12544 18629 13568
rect 18309 12480 18317 12544
rect 18381 12480 18397 12544
rect 18461 12480 18477 12544
rect 18541 12480 18557 12544
rect 18621 12480 18629 12544
rect 18309 11456 18629 12480
rect 18309 11392 18317 11456
rect 18381 11392 18397 11456
rect 18461 11392 18477 11456
rect 18541 11392 18557 11456
rect 18621 11392 18629 11456
rect 18309 10368 18629 11392
rect 18309 10304 18317 10368
rect 18381 10304 18397 10368
rect 18461 10304 18477 10368
rect 18541 10304 18557 10368
rect 18621 10304 18629 10368
rect 18309 9280 18629 10304
rect 18309 9216 18317 9280
rect 18381 9216 18397 9280
rect 18461 9216 18477 9280
rect 18541 9216 18557 9280
rect 18621 9216 18629 9280
rect 18309 8192 18629 9216
rect 18309 8128 18317 8192
rect 18381 8128 18397 8192
rect 18461 8128 18477 8192
rect 18541 8128 18557 8192
rect 18621 8128 18629 8192
rect 18309 7104 18629 8128
rect 18309 7040 18317 7104
rect 18381 7040 18397 7104
rect 18461 7040 18477 7104
rect 18541 7040 18557 7104
rect 18621 7040 18629 7104
rect 18309 6016 18629 7040
rect 18309 5952 18317 6016
rect 18381 5952 18397 6016
rect 18461 5952 18477 6016
rect 18541 5952 18557 6016
rect 18621 5952 18629 6016
rect 18309 4928 18629 5952
rect 18309 4864 18317 4928
rect 18381 4864 18397 4928
rect 18461 4864 18477 4928
rect 18541 4864 18557 4928
rect 18621 4864 18629 4928
rect 18309 3840 18629 4864
rect 18309 3776 18317 3840
rect 18381 3776 18397 3840
rect 18461 3776 18477 3840
rect 18541 3776 18557 3840
rect 18621 3776 18629 3840
rect 18309 2752 18629 3776
rect 18309 2688 18317 2752
rect 18381 2688 18397 2752
rect 18461 2688 18477 2752
rect 18541 2688 18557 2752
rect 18621 2688 18629 2752
rect 18309 2128 18629 2688
rect 21782 31584 22102 31600
rect 21782 31520 21790 31584
rect 21854 31520 21870 31584
rect 21934 31520 21950 31584
rect 22014 31520 22030 31584
rect 22094 31520 22102 31584
rect 21782 30496 22102 31520
rect 21782 30432 21790 30496
rect 21854 30432 21870 30496
rect 21934 30432 21950 30496
rect 22014 30432 22030 30496
rect 22094 30432 22102 30496
rect 21782 29408 22102 30432
rect 21782 29344 21790 29408
rect 21854 29344 21870 29408
rect 21934 29344 21950 29408
rect 22014 29344 22030 29408
rect 22094 29344 22102 29408
rect 21782 28320 22102 29344
rect 21782 28256 21790 28320
rect 21854 28256 21870 28320
rect 21934 28256 21950 28320
rect 22014 28256 22030 28320
rect 22094 28256 22102 28320
rect 21782 27232 22102 28256
rect 21782 27168 21790 27232
rect 21854 27168 21870 27232
rect 21934 27168 21950 27232
rect 22014 27168 22030 27232
rect 22094 27168 22102 27232
rect 21782 26144 22102 27168
rect 21782 26080 21790 26144
rect 21854 26080 21870 26144
rect 21934 26080 21950 26144
rect 22014 26080 22030 26144
rect 22094 26080 22102 26144
rect 21782 25056 22102 26080
rect 21782 24992 21790 25056
rect 21854 24992 21870 25056
rect 21934 24992 21950 25056
rect 22014 24992 22030 25056
rect 22094 24992 22102 25056
rect 21782 23968 22102 24992
rect 21782 23904 21790 23968
rect 21854 23904 21870 23968
rect 21934 23904 21950 23968
rect 22014 23904 22030 23968
rect 22094 23904 22102 23968
rect 21782 22880 22102 23904
rect 21782 22816 21790 22880
rect 21854 22816 21870 22880
rect 21934 22816 21950 22880
rect 22014 22816 22030 22880
rect 22094 22816 22102 22880
rect 21782 21792 22102 22816
rect 21782 21728 21790 21792
rect 21854 21728 21870 21792
rect 21934 21728 21950 21792
rect 22014 21728 22030 21792
rect 22094 21728 22102 21792
rect 21782 20704 22102 21728
rect 21782 20640 21790 20704
rect 21854 20640 21870 20704
rect 21934 20640 21950 20704
rect 22014 20640 22030 20704
rect 22094 20640 22102 20704
rect 21782 19616 22102 20640
rect 21782 19552 21790 19616
rect 21854 19552 21870 19616
rect 21934 19552 21950 19616
rect 22014 19552 22030 19616
rect 22094 19552 22102 19616
rect 21782 18528 22102 19552
rect 21782 18464 21790 18528
rect 21854 18464 21870 18528
rect 21934 18464 21950 18528
rect 22014 18464 22030 18528
rect 22094 18464 22102 18528
rect 21782 17440 22102 18464
rect 21782 17376 21790 17440
rect 21854 17376 21870 17440
rect 21934 17376 21950 17440
rect 22014 17376 22030 17440
rect 22094 17376 22102 17440
rect 21782 16352 22102 17376
rect 21782 16288 21790 16352
rect 21854 16288 21870 16352
rect 21934 16288 21950 16352
rect 22014 16288 22030 16352
rect 22094 16288 22102 16352
rect 21782 15264 22102 16288
rect 21782 15200 21790 15264
rect 21854 15200 21870 15264
rect 21934 15200 21950 15264
rect 22014 15200 22030 15264
rect 22094 15200 22102 15264
rect 21782 14176 22102 15200
rect 21782 14112 21790 14176
rect 21854 14112 21870 14176
rect 21934 14112 21950 14176
rect 22014 14112 22030 14176
rect 22094 14112 22102 14176
rect 21782 13088 22102 14112
rect 21782 13024 21790 13088
rect 21854 13024 21870 13088
rect 21934 13024 21950 13088
rect 22014 13024 22030 13088
rect 22094 13024 22102 13088
rect 21782 12000 22102 13024
rect 21782 11936 21790 12000
rect 21854 11936 21870 12000
rect 21934 11936 21950 12000
rect 22014 11936 22030 12000
rect 22094 11936 22102 12000
rect 21782 10912 22102 11936
rect 21782 10848 21790 10912
rect 21854 10848 21870 10912
rect 21934 10848 21950 10912
rect 22014 10848 22030 10912
rect 22094 10848 22102 10912
rect 21782 9824 22102 10848
rect 21782 9760 21790 9824
rect 21854 9760 21870 9824
rect 21934 9760 21950 9824
rect 22014 9760 22030 9824
rect 22094 9760 22102 9824
rect 21782 8736 22102 9760
rect 21782 8672 21790 8736
rect 21854 8672 21870 8736
rect 21934 8672 21950 8736
rect 22014 8672 22030 8736
rect 22094 8672 22102 8736
rect 21782 7648 22102 8672
rect 21782 7584 21790 7648
rect 21854 7584 21870 7648
rect 21934 7584 21950 7648
rect 22014 7584 22030 7648
rect 22094 7584 22102 7648
rect 21782 6560 22102 7584
rect 21782 6496 21790 6560
rect 21854 6496 21870 6560
rect 21934 6496 21950 6560
rect 22014 6496 22030 6560
rect 22094 6496 22102 6560
rect 21782 5472 22102 6496
rect 21782 5408 21790 5472
rect 21854 5408 21870 5472
rect 21934 5408 21950 5472
rect 22014 5408 22030 5472
rect 22094 5408 22102 5472
rect 21782 4384 22102 5408
rect 21782 4320 21790 4384
rect 21854 4320 21870 4384
rect 21934 4320 21950 4384
rect 22014 4320 22030 4384
rect 22094 4320 22102 4384
rect 21782 3296 22102 4320
rect 21782 3232 21790 3296
rect 21854 3232 21870 3296
rect 21934 3232 21950 3296
rect 22014 3232 22030 3296
rect 22094 3232 22102 3296
rect 21782 2208 22102 3232
rect 21782 2144 21790 2208
rect 21854 2144 21870 2208
rect 21934 2144 21950 2208
rect 22014 2144 22030 2208
rect 22094 2144 22102 2208
rect 21782 2128 22102 2144
rect 25255 31040 25575 31600
rect 25255 30976 25263 31040
rect 25327 30976 25343 31040
rect 25407 30976 25423 31040
rect 25487 30976 25503 31040
rect 25567 30976 25575 31040
rect 25255 29952 25575 30976
rect 25255 29888 25263 29952
rect 25327 29888 25343 29952
rect 25407 29888 25423 29952
rect 25487 29888 25503 29952
rect 25567 29888 25575 29952
rect 25255 28864 25575 29888
rect 25255 28800 25263 28864
rect 25327 28800 25343 28864
rect 25407 28800 25423 28864
rect 25487 28800 25503 28864
rect 25567 28800 25575 28864
rect 25255 27776 25575 28800
rect 25255 27712 25263 27776
rect 25327 27712 25343 27776
rect 25407 27712 25423 27776
rect 25487 27712 25503 27776
rect 25567 27712 25575 27776
rect 25255 26688 25575 27712
rect 25255 26624 25263 26688
rect 25327 26624 25343 26688
rect 25407 26624 25423 26688
rect 25487 26624 25503 26688
rect 25567 26624 25575 26688
rect 25255 25600 25575 26624
rect 25255 25536 25263 25600
rect 25327 25536 25343 25600
rect 25407 25536 25423 25600
rect 25487 25536 25503 25600
rect 25567 25536 25575 25600
rect 25255 24512 25575 25536
rect 25255 24448 25263 24512
rect 25327 24448 25343 24512
rect 25407 24448 25423 24512
rect 25487 24448 25503 24512
rect 25567 24448 25575 24512
rect 25255 23424 25575 24448
rect 25255 23360 25263 23424
rect 25327 23360 25343 23424
rect 25407 23360 25423 23424
rect 25487 23360 25503 23424
rect 25567 23360 25575 23424
rect 25255 22336 25575 23360
rect 25255 22272 25263 22336
rect 25327 22272 25343 22336
rect 25407 22272 25423 22336
rect 25487 22272 25503 22336
rect 25567 22272 25575 22336
rect 25255 21248 25575 22272
rect 25255 21184 25263 21248
rect 25327 21184 25343 21248
rect 25407 21184 25423 21248
rect 25487 21184 25503 21248
rect 25567 21184 25575 21248
rect 25255 20160 25575 21184
rect 25255 20096 25263 20160
rect 25327 20096 25343 20160
rect 25407 20096 25423 20160
rect 25487 20096 25503 20160
rect 25567 20096 25575 20160
rect 25255 19072 25575 20096
rect 25255 19008 25263 19072
rect 25327 19008 25343 19072
rect 25407 19008 25423 19072
rect 25487 19008 25503 19072
rect 25567 19008 25575 19072
rect 25255 17984 25575 19008
rect 25255 17920 25263 17984
rect 25327 17920 25343 17984
rect 25407 17920 25423 17984
rect 25487 17920 25503 17984
rect 25567 17920 25575 17984
rect 25255 16896 25575 17920
rect 25255 16832 25263 16896
rect 25327 16832 25343 16896
rect 25407 16832 25423 16896
rect 25487 16832 25503 16896
rect 25567 16832 25575 16896
rect 25255 15808 25575 16832
rect 25255 15744 25263 15808
rect 25327 15744 25343 15808
rect 25407 15744 25423 15808
rect 25487 15744 25503 15808
rect 25567 15744 25575 15808
rect 25255 14720 25575 15744
rect 25255 14656 25263 14720
rect 25327 14656 25343 14720
rect 25407 14656 25423 14720
rect 25487 14656 25503 14720
rect 25567 14656 25575 14720
rect 25255 13632 25575 14656
rect 25255 13568 25263 13632
rect 25327 13568 25343 13632
rect 25407 13568 25423 13632
rect 25487 13568 25503 13632
rect 25567 13568 25575 13632
rect 25255 12544 25575 13568
rect 25255 12480 25263 12544
rect 25327 12480 25343 12544
rect 25407 12480 25423 12544
rect 25487 12480 25503 12544
rect 25567 12480 25575 12544
rect 25255 11456 25575 12480
rect 25255 11392 25263 11456
rect 25327 11392 25343 11456
rect 25407 11392 25423 11456
rect 25487 11392 25503 11456
rect 25567 11392 25575 11456
rect 25255 10368 25575 11392
rect 25255 10304 25263 10368
rect 25327 10304 25343 10368
rect 25407 10304 25423 10368
rect 25487 10304 25503 10368
rect 25567 10304 25575 10368
rect 25255 9280 25575 10304
rect 25255 9216 25263 9280
rect 25327 9216 25343 9280
rect 25407 9216 25423 9280
rect 25487 9216 25503 9280
rect 25567 9216 25575 9280
rect 25255 8192 25575 9216
rect 25255 8128 25263 8192
rect 25327 8128 25343 8192
rect 25407 8128 25423 8192
rect 25487 8128 25503 8192
rect 25567 8128 25575 8192
rect 25255 7104 25575 8128
rect 25255 7040 25263 7104
rect 25327 7040 25343 7104
rect 25407 7040 25423 7104
rect 25487 7040 25503 7104
rect 25567 7040 25575 7104
rect 25255 6016 25575 7040
rect 25255 5952 25263 6016
rect 25327 5952 25343 6016
rect 25407 5952 25423 6016
rect 25487 5952 25503 6016
rect 25567 5952 25575 6016
rect 25255 4928 25575 5952
rect 25255 4864 25263 4928
rect 25327 4864 25343 4928
rect 25407 4864 25423 4928
rect 25487 4864 25503 4928
rect 25567 4864 25575 4928
rect 25255 3840 25575 4864
rect 25255 3776 25263 3840
rect 25327 3776 25343 3840
rect 25407 3776 25423 3840
rect 25487 3776 25503 3840
rect 25567 3776 25575 3840
rect 25255 2752 25575 3776
rect 25255 2688 25263 2752
rect 25327 2688 25343 2752
rect 25407 2688 25423 2752
rect 25487 2688 25503 2752
rect 25567 2688 25575 2752
rect 25255 2128 25575 2688
rect 28728 31584 29048 31600
rect 28728 31520 28736 31584
rect 28800 31520 28816 31584
rect 28880 31520 28896 31584
rect 28960 31520 28976 31584
rect 29040 31520 29048 31584
rect 28728 30496 29048 31520
rect 28728 30432 28736 30496
rect 28800 30432 28816 30496
rect 28880 30432 28896 30496
rect 28960 30432 28976 30496
rect 29040 30432 29048 30496
rect 28728 29408 29048 30432
rect 28728 29344 28736 29408
rect 28800 29344 28816 29408
rect 28880 29344 28896 29408
rect 28960 29344 28976 29408
rect 29040 29344 29048 29408
rect 28728 28320 29048 29344
rect 28728 28256 28736 28320
rect 28800 28256 28816 28320
rect 28880 28256 28896 28320
rect 28960 28256 28976 28320
rect 29040 28256 29048 28320
rect 28728 27232 29048 28256
rect 28728 27168 28736 27232
rect 28800 27168 28816 27232
rect 28880 27168 28896 27232
rect 28960 27168 28976 27232
rect 29040 27168 29048 27232
rect 28728 26144 29048 27168
rect 28728 26080 28736 26144
rect 28800 26080 28816 26144
rect 28880 26080 28896 26144
rect 28960 26080 28976 26144
rect 29040 26080 29048 26144
rect 28728 25056 29048 26080
rect 28728 24992 28736 25056
rect 28800 24992 28816 25056
rect 28880 24992 28896 25056
rect 28960 24992 28976 25056
rect 29040 24992 29048 25056
rect 28728 23968 29048 24992
rect 28728 23904 28736 23968
rect 28800 23904 28816 23968
rect 28880 23904 28896 23968
rect 28960 23904 28976 23968
rect 29040 23904 29048 23968
rect 28728 22880 29048 23904
rect 28728 22816 28736 22880
rect 28800 22816 28816 22880
rect 28880 22816 28896 22880
rect 28960 22816 28976 22880
rect 29040 22816 29048 22880
rect 28728 21792 29048 22816
rect 28728 21728 28736 21792
rect 28800 21728 28816 21792
rect 28880 21728 28896 21792
rect 28960 21728 28976 21792
rect 29040 21728 29048 21792
rect 28728 20704 29048 21728
rect 28728 20640 28736 20704
rect 28800 20640 28816 20704
rect 28880 20640 28896 20704
rect 28960 20640 28976 20704
rect 29040 20640 29048 20704
rect 28728 19616 29048 20640
rect 28728 19552 28736 19616
rect 28800 19552 28816 19616
rect 28880 19552 28896 19616
rect 28960 19552 28976 19616
rect 29040 19552 29048 19616
rect 28728 18528 29048 19552
rect 28728 18464 28736 18528
rect 28800 18464 28816 18528
rect 28880 18464 28896 18528
rect 28960 18464 28976 18528
rect 29040 18464 29048 18528
rect 28728 17440 29048 18464
rect 28728 17376 28736 17440
rect 28800 17376 28816 17440
rect 28880 17376 28896 17440
rect 28960 17376 28976 17440
rect 29040 17376 29048 17440
rect 28728 16352 29048 17376
rect 28728 16288 28736 16352
rect 28800 16288 28816 16352
rect 28880 16288 28896 16352
rect 28960 16288 28976 16352
rect 29040 16288 29048 16352
rect 28728 15264 29048 16288
rect 28728 15200 28736 15264
rect 28800 15200 28816 15264
rect 28880 15200 28896 15264
rect 28960 15200 28976 15264
rect 29040 15200 29048 15264
rect 28728 14176 29048 15200
rect 28728 14112 28736 14176
rect 28800 14112 28816 14176
rect 28880 14112 28896 14176
rect 28960 14112 28976 14176
rect 29040 14112 29048 14176
rect 28728 13088 29048 14112
rect 28728 13024 28736 13088
rect 28800 13024 28816 13088
rect 28880 13024 28896 13088
rect 28960 13024 28976 13088
rect 29040 13024 29048 13088
rect 28728 12000 29048 13024
rect 28728 11936 28736 12000
rect 28800 11936 28816 12000
rect 28880 11936 28896 12000
rect 28960 11936 28976 12000
rect 29040 11936 29048 12000
rect 28728 10912 29048 11936
rect 28728 10848 28736 10912
rect 28800 10848 28816 10912
rect 28880 10848 28896 10912
rect 28960 10848 28976 10912
rect 29040 10848 29048 10912
rect 28728 9824 29048 10848
rect 28728 9760 28736 9824
rect 28800 9760 28816 9824
rect 28880 9760 28896 9824
rect 28960 9760 28976 9824
rect 29040 9760 29048 9824
rect 28728 8736 29048 9760
rect 28728 8672 28736 8736
rect 28800 8672 28816 8736
rect 28880 8672 28896 8736
rect 28960 8672 28976 8736
rect 29040 8672 29048 8736
rect 28728 7648 29048 8672
rect 28728 7584 28736 7648
rect 28800 7584 28816 7648
rect 28880 7584 28896 7648
rect 28960 7584 28976 7648
rect 29040 7584 29048 7648
rect 28728 6560 29048 7584
rect 28728 6496 28736 6560
rect 28800 6496 28816 6560
rect 28880 6496 28896 6560
rect 28960 6496 28976 6560
rect 29040 6496 29048 6560
rect 28728 5472 29048 6496
rect 28728 5408 28736 5472
rect 28800 5408 28816 5472
rect 28880 5408 28896 5472
rect 28960 5408 28976 5472
rect 29040 5408 29048 5472
rect 28728 4384 29048 5408
rect 28728 4320 28736 4384
rect 28800 4320 28816 4384
rect 28880 4320 28896 4384
rect 28960 4320 28976 4384
rect 29040 4320 29048 4384
rect 28728 3296 29048 4320
rect 28728 3232 28736 3296
rect 28800 3232 28816 3296
rect 28880 3232 28896 3296
rect 28960 3232 28976 3296
rect 29040 3232 29048 3296
rect 28728 2208 29048 3232
rect 28728 2144 28736 2208
rect 28800 2144 28816 2208
rect 28880 2144 28896 2208
rect 28960 2144 28976 2208
rect 29040 2144 29048 2208
rect 28728 2128 29048 2144
rect 12755 1460 12821 1461
rect 12755 1396 12756 1460
rect 12820 1396 12821 1460
rect 12755 1395 12821 1396
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 17572 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1666464484
transform -1 0 4416 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__B
timestamp 1666464484
transform 1 0 15456 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1666464484
transform 1 0 4784 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__B1
timestamp 1666464484
transform 1 0 13616 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1666464484
transform 1 0 13248 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1666464484
transform 1 0 13248 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1666464484
transform 1 0 11040 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__B
timestamp 1666464484
transform 1 0 13524 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1666464484
transform 1 0 12420 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__B
timestamp 1666464484
transform -1 0 12328 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A1
timestamp 1666464484
transform -1 0 11408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A2
timestamp 1666464484
transform 1 0 10028 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__B1
timestamp 1666464484
transform -1 0 11132 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__B
timestamp 1666464484
transform -1 0 20700 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__C
timestamp 1666464484
transform -1 0 21528 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1666464484
transform -1 0 20700 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1666464484
transform -1 0 18400 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1666464484
transform 1 0 18216 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A1
timestamp 1666464484
transform 1 0 11132 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__B
timestamp 1666464484
transform 1 0 10948 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__B
timestamp 1666464484
transform 1 0 5152 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__C
timestamp 1666464484
transform -1 0 5152 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__B1
timestamp 1666464484
transform 1 0 6532 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A
timestamp 1666464484
transform -1 0 10580 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A2
timestamp 1666464484
transform -1 0 17480 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__B1
timestamp 1666464484
transform 1 0 16192 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__A2
timestamp 1666464484
transform 1 0 2392 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A2
timestamp 1666464484
transform 1 0 3864 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__C
timestamp 1666464484
transform 1 0 14260 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1666464484
transform 1 0 5428 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__B1
timestamp 1666464484
transform 1 0 14628 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__130__C
timestamp 1666464484
transform 1 0 11684 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__131__A
timestamp 1666464484
transform 1 0 4416 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__133__B1
timestamp 1666464484
transform -1 0 17020 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__136__A
timestamp 1666464484
transform 1 0 17664 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__A
timestamp 1666464484
transform 1 0 19964 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__B1
timestamp 1666464484
transform -1 0 9384 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__145__A
timestamp 1666464484
transform 1 0 14904 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__149__A
timestamp 1666464484
transform 1 0 4232 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__B1
timestamp 1666464484
transform -1 0 6532 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__A
timestamp 1666464484
transform 1 0 3312 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__C
timestamp 1666464484
transform -1 0 3496 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__A
timestamp 1666464484
transform 1 0 14076 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__A2
timestamp 1666464484
transform -1 0 20148 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__160__B1
timestamp 1666464484
transform 1 0 19412 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__164__A
timestamp 1666464484
transform -1 0 20976 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__167__A
timestamp 1666464484
transform -1 0 6992 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__169__B1
timestamp 1666464484
transform 1 0 2576 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__A
timestamp 1666464484
transform 1 0 5888 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__176__A
timestamp 1666464484
transform -1 0 8832 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__179__A
timestamp 1666464484
transform 1 0 6992 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__A1
timestamp 1666464484
transform 1 0 9108 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__B1
timestamp 1666464484
transform -1 0 7912 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__182__A1
timestamp 1666464484
transform -1 0 2208 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__183__A1
timestamp 1666464484
transform -1 0 9660 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__A2
timestamp 1666464484
transform 1 0 8464 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__B1
timestamp 1666464484
transform 1 0 10028 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__186__D
timestamp 1666464484
transform 1 0 4232 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__D
timestamp 1666464484
transform 1 0 11132 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_io_in[0]_A
timestamp 1666464484
transform -1 0 11224 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1666464484
transform -1 0 28428 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1666464484
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1666464484
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1666464484
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1666464484
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1666464484
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1666464484
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1666464484
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1666464484
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1666464484
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1666464484
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1666464484
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1666464484
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1666464484
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1666464484
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1666464484
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1666464484
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1666464484
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1666464484
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1666464484
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1666464484
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1666464484
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1666464484
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1666464484
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1666464484
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1666464484
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1666464484
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1666464484
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1666464484
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_293 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28060 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1666464484
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1666464484
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1666464484
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1666464484
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1666464484
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1666464484
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1666464484
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1666464484
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1666464484
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1666464484
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1666464484
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1666464484
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1666464484
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1666464484
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1666464484
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1666464484
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1666464484
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1666464484
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1666464484
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1666464484
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1666464484
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1666464484
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1666464484
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1666464484
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1666464484
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1666464484
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1666464484
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1666464484
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1666464484
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1666464484
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_293
timestamp 1666464484
transform 1 0 28060 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_297 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28428 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1666464484
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_8
timestamp 1666464484
transform 1 0 1840 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1666464484
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1666464484
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1666464484
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1666464484
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1666464484
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1666464484
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1666464484
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1666464484
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1666464484
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1666464484
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1666464484
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1666464484
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1666464484
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1666464484
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1666464484
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1666464484
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1666464484
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1666464484
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1666464484
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1666464484
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1666464484
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1666464484
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1666464484
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1666464484
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1666464484
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1666464484
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1666464484
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_289
timestamp 1666464484
transform 1 0 27692 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_293
timestamp 1666464484
transform 1 0 28060 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_297
timestamp 1666464484
transform 1 0 28428 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1666464484
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_8
timestamp 1666464484
transform 1 0 1840 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_20
timestamp 1666464484
transform 1 0 2944 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_32
timestamp 1666464484
transform 1 0 4048 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_44
timestamp 1666464484
transform 1 0 5152 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1666464484
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1666464484
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1666464484
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1666464484
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1666464484
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1666464484
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1666464484
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1666464484
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1666464484
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1666464484
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1666464484
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1666464484
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1666464484
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1666464484
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1666464484
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1666464484
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1666464484
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1666464484
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1666464484
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1666464484
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1666464484
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1666464484
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1666464484
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1666464484
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_281
timestamp 1666464484
transform 1 0 26956 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_297
timestamp 1666464484
transform 1 0 28428 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1666464484
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1666464484
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1666464484
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1666464484
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1666464484
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1666464484
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1666464484
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1666464484
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1666464484
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1666464484
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1666464484
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1666464484
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1666464484
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1666464484
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1666464484
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1666464484
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1666464484
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1666464484
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1666464484
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1666464484
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1666464484
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1666464484
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1666464484
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1666464484
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1666464484
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1666464484
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1666464484
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1666464484
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1666464484
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1666464484
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_289
timestamp 1666464484
transform 1 0 27692 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_297
timestamp 1666464484
transform 1 0 28428 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1666464484
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_8
timestamp 1666464484
transform 1 0 1840 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_20
timestamp 1666464484
transform 1 0 2944 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_32
timestamp 1666464484
transform 1 0 4048 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_44
timestamp 1666464484
transform 1 0 5152 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1666464484
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1666464484
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1666464484
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1666464484
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1666464484
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1666464484
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1666464484
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1666464484
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1666464484
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1666464484
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1666464484
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1666464484
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1666464484
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1666464484
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1666464484
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1666464484
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1666464484
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1666464484
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1666464484
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1666464484
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1666464484
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1666464484
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1666464484
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1666464484
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1666464484
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_293
timestamp 1666464484
transform 1 0 28060 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_297
timestamp 1666464484
transform 1 0 28428 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1666464484
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1666464484
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1666464484
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1666464484
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1666464484
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1666464484
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1666464484
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1666464484
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1666464484
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1666464484
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1666464484
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1666464484
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1666464484
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1666464484
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1666464484
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1666464484
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1666464484
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1666464484
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1666464484
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1666464484
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1666464484
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1666464484
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1666464484
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1666464484
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1666464484
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1666464484
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1666464484
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1666464484
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1666464484
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1666464484
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_289
timestamp 1666464484
transform 1 0 27692 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_293
timestamp 1666464484
transform 1 0 28060 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_297
timestamp 1666464484
transform 1 0 28428 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1666464484
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_8
timestamp 1666464484
transform 1 0 1840 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_20
timestamp 1666464484
transform 1 0 2944 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_32
timestamp 1666464484
transform 1 0 4048 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_44
timestamp 1666464484
transform 1 0 5152 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1666464484
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1666464484
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1666464484
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1666464484
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1666464484
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1666464484
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1666464484
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1666464484
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1666464484
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1666464484
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1666464484
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1666464484
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1666464484
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1666464484
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1666464484
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1666464484
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1666464484
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1666464484
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1666464484
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1666464484
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1666464484
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1666464484
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1666464484
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1666464484
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1666464484
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_293
timestamp 1666464484
transform 1 0 28060 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1666464484
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1666464484
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1666464484
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1666464484
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1666464484
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1666464484
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1666464484
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1666464484
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1666464484
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1666464484
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1666464484
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1666464484
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1666464484
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1666464484
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1666464484
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1666464484
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1666464484
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1666464484
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1666464484
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1666464484
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1666464484
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1666464484
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1666464484
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1666464484
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1666464484
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1666464484
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1666464484
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1666464484
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1666464484
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1666464484
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_289
timestamp 1666464484
transform 1 0 27692 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_293
timestamp 1666464484
transform 1 0 28060 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_297
timestamp 1666464484
transform 1 0 28428 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1666464484
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_8
timestamp 1666464484
transform 1 0 1840 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_20
timestamp 1666464484
transform 1 0 2944 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_32
timestamp 1666464484
transform 1 0 4048 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_44
timestamp 1666464484
transform 1 0 5152 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1666464484
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1666464484
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1666464484
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1666464484
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1666464484
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1666464484
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1666464484
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1666464484
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1666464484
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1666464484
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1666464484
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1666464484
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1666464484
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1666464484
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1666464484
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1666464484
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1666464484
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1666464484
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1666464484
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1666464484
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1666464484
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1666464484
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1666464484
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1666464484
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1666464484
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_293
timestamp 1666464484
transform 1 0 28060 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1666464484
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_8
timestamp 1666464484
transform 1 0 1840 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_20
timestamp 1666464484
transform 1 0 2944 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1666464484
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1666464484
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1666464484
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1666464484
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1666464484
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1666464484
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1666464484
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1666464484
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1666464484
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1666464484
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1666464484
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1666464484
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1666464484
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1666464484
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1666464484
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1666464484
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1666464484
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1666464484
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1666464484
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1666464484
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1666464484
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1666464484
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1666464484
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1666464484
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1666464484
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1666464484
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1666464484
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_289
timestamp 1666464484
transform 1 0 27692 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_293
timestamp 1666464484
transform 1 0 28060 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_297
timestamp 1666464484
transform 1 0 28428 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1666464484
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1666464484
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1666464484
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1666464484
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1666464484
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1666464484
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1666464484
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1666464484
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1666464484
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1666464484
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1666464484
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1666464484
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1666464484
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1666464484
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1666464484
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1666464484
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1666464484
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1666464484
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1666464484
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1666464484
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1666464484
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1666464484
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1666464484
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1666464484
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1666464484
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1666464484
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1666464484
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1666464484
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1666464484
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1666464484
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1666464484
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_293
timestamp 1666464484
transform 1 0 28060 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1666464484
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1666464484
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1666464484
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1666464484
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1666464484
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1666464484
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1666464484
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1666464484
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1666464484
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1666464484
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1666464484
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1666464484
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1666464484
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1666464484
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1666464484
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1666464484
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1666464484
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1666464484
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1666464484
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1666464484
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1666464484
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1666464484
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1666464484
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1666464484
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1666464484
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1666464484
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1666464484
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1666464484
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1666464484
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1666464484
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_289
timestamp 1666464484
transform 1 0 27692 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_293
timestamp 1666464484
transform 1 0 28060 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_297
timestamp 1666464484
transform 1 0 28428 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1666464484
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_8
timestamp 1666464484
transform 1 0 1840 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_20
timestamp 1666464484
transform 1 0 2944 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_32
timestamp 1666464484
transform 1 0 4048 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_44
timestamp 1666464484
transform 1 0 5152 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1666464484
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1666464484
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1666464484
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1666464484
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1666464484
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1666464484
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1666464484
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1666464484
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1666464484
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1666464484
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1666464484
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1666464484
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1666464484
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1666464484
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1666464484
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1666464484
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1666464484
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1666464484
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1666464484
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1666464484
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1666464484
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1666464484
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1666464484
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1666464484
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1666464484
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_293
timestamp 1666464484
transform 1 0 28060 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_297
timestamp 1666464484
transform 1 0 28428 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1666464484
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_8
timestamp 1666464484
transform 1 0 1840 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_20
timestamp 1666464484
transform 1 0 2944 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1666464484
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1666464484
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1666464484
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1666464484
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1666464484
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1666464484
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1666464484
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1666464484
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1666464484
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1666464484
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1666464484
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1666464484
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1666464484
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1666464484
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1666464484
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1666464484
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1666464484
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1666464484
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1666464484
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1666464484
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1666464484
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1666464484
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1666464484
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1666464484
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1666464484
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1666464484
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1666464484
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_289
timestamp 1666464484
transform 1 0 27692 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_297
timestamp 1666464484
transform 1 0 28428 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1666464484
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1666464484
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1666464484
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1666464484
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1666464484
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1666464484
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1666464484
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1666464484
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1666464484
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1666464484
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1666464484
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1666464484
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1666464484
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1666464484
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1666464484
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1666464484
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1666464484
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1666464484
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1666464484
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1666464484
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1666464484
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1666464484
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1666464484
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1666464484
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1666464484
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1666464484
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1666464484
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1666464484
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1666464484
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1666464484
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1666464484
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_293
timestamp 1666464484
transform 1 0 28060 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1666464484
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1666464484
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1666464484
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1666464484
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1666464484
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1666464484
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1666464484
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1666464484
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1666464484
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1666464484
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1666464484
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1666464484
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1666464484
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1666464484
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1666464484
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1666464484
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1666464484
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1666464484
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1666464484
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1666464484
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1666464484
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1666464484
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1666464484
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1666464484
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1666464484
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1666464484
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1666464484
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1666464484
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1666464484
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1666464484
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_289
timestamp 1666464484
transform 1 0 27692 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_293
timestamp 1666464484
transform 1 0 28060 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_297
timestamp 1666464484
transform 1 0 28428 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1666464484
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_8
timestamp 1666464484
transform 1 0 1840 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_20
timestamp 1666464484
transform 1 0 2944 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_32
timestamp 1666464484
transform 1 0 4048 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_44
timestamp 1666464484
transform 1 0 5152 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1666464484
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1666464484
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1666464484
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1666464484
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1666464484
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1666464484
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1666464484
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1666464484
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1666464484
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1666464484
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1666464484
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1666464484
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1666464484
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1666464484
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1666464484
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1666464484
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1666464484
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1666464484
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1666464484
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1666464484
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1666464484
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1666464484
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1666464484
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1666464484
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1666464484
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_293
timestamp 1666464484
transform 1 0 28060 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_297
timestamp 1666464484
transform 1 0 28428 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1666464484
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_8
timestamp 1666464484
transform 1 0 1840 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_20
timestamp 1666464484
transform 1 0 2944 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1666464484
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1666464484
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1666464484
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1666464484
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1666464484
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1666464484
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1666464484
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1666464484
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1666464484
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1666464484
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1666464484
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1666464484
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1666464484
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1666464484
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1666464484
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1666464484
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1666464484
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1666464484
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1666464484
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1666464484
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1666464484
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1666464484
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1666464484
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1666464484
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1666464484
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1666464484
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1666464484
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_289
timestamp 1666464484
transform 1 0 27692 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_297
timestamp 1666464484
transform 1 0 28428 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1666464484
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1666464484
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1666464484
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1666464484
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1666464484
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1666464484
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1666464484
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1666464484
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1666464484
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1666464484
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1666464484
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1666464484
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1666464484
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1666464484
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1666464484
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1666464484
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1666464484
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1666464484
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1666464484
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1666464484
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1666464484
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1666464484
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1666464484
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1666464484
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1666464484
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1666464484
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1666464484
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1666464484
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1666464484
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1666464484
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1666464484
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_293
timestamp 1666464484
transform 1 0 28060 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1666464484
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_8
timestamp 1666464484
transform 1 0 1840 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_20
timestamp 1666464484
transform 1 0 2944 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1666464484
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1666464484
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1666464484
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1666464484
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1666464484
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1666464484
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1666464484
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1666464484
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1666464484
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1666464484
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1666464484
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1666464484
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1666464484
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1666464484
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1666464484
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1666464484
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1666464484
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1666464484
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1666464484
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1666464484
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1666464484
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1666464484
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1666464484
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1666464484
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1666464484
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1666464484
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1666464484
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_289
timestamp 1666464484
transform 1 0 27692 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_293
timestamp 1666464484
transform 1 0 28060 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_297
timestamp 1666464484
transform 1 0 28428 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1666464484
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1666464484
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1666464484
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1666464484
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1666464484
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1666464484
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1666464484
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1666464484
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1666464484
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1666464484
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1666464484
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1666464484
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1666464484
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1666464484
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1666464484
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1666464484
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1666464484
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1666464484
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1666464484
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1666464484
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1666464484
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1666464484
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1666464484
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1666464484
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1666464484
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1666464484
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1666464484
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1666464484
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1666464484
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1666464484
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1666464484
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_293
timestamp 1666464484
transform 1 0 28060 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_297
timestamp 1666464484
transform 1 0 28428 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1666464484
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_8
timestamp 1666464484
transform 1 0 1840 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_20
timestamp 1666464484
transform 1 0 2944 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1666464484
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1666464484
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1666464484
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1666464484
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1666464484
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1666464484
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1666464484
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1666464484
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1666464484
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1666464484
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1666464484
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1666464484
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1666464484
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1666464484
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1666464484
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1666464484
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1666464484
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1666464484
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1666464484
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1666464484
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1666464484
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1666464484
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1666464484
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1666464484
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1666464484
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1666464484
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1666464484
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_289
timestamp 1666464484
transform 1 0 27692 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_297
timestamp 1666464484
transform 1 0 28428 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1666464484
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1666464484
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1666464484
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1666464484
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1666464484
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1666464484
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1666464484
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1666464484
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1666464484
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1666464484
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1666464484
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1666464484
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1666464484
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1666464484
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1666464484
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1666464484
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1666464484
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1666464484
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1666464484
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1666464484
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1666464484
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1666464484
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1666464484
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1666464484
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1666464484
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1666464484
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1666464484
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1666464484
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1666464484
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1666464484
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1666464484
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_293
timestamp 1666464484
transform 1 0 28060 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_297
timestamp 1666464484
transform 1 0 28428 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1666464484
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_8
timestamp 1666464484
transform 1 0 1840 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_20
timestamp 1666464484
transform 1 0 2944 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1666464484
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1666464484
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1666464484
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1666464484
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1666464484
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1666464484
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1666464484
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1666464484
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1666464484
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1666464484
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1666464484
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1666464484
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1666464484
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1666464484
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1666464484
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1666464484
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1666464484
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1666464484
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1666464484
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1666464484
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1666464484
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1666464484
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1666464484
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1666464484
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1666464484
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1666464484
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1666464484
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_289
timestamp 1666464484
transform 1 0 27692 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_297
timestamp 1666464484
transform 1 0 28428 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1666464484
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_8
timestamp 1666464484
transform 1 0 1840 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_20
timestamp 1666464484
transform 1 0 2944 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_32
timestamp 1666464484
transform 1 0 4048 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_44
timestamp 1666464484
transform 1 0 5152 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1666464484
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1666464484
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1666464484
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1666464484
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1666464484
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1666464484
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1666464484
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1666464484
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1666464484
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1666464484
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1666464484
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1666464484
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1666464484
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1666464484
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1666464484
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1666464484
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1666464484
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1666464484
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1666464484
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1666464484
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1666464484
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1666464484
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1666464484
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1666464484
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1666464484
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_293
timestamp 1666464484
transform 1 0 28060 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_297
timestamp 1666464484
transform 1 0 28428 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1666464484
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1666464484
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1666464484
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1666464484
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1666464484
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1666464484
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1666464484
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1666464484
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1666464484
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1666464484
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1666464484
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1666464484
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1666464484
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1666464484
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1666464484
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1666464484
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1666464484
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1666464484
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1666464484
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1666464484
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1666464484
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1666464484
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1666464484
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1666464484
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1666464484
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1666464484
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1666464484
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1666464484
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1666464484
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1666464484
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_289
timestamp 1666464484
transform 1 0 27692 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_297
timestamp 1666464484
transform 1 0 28428 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1666464484
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1666464484
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1666464484
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1666464484
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1666464484
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1666464484
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1666464484
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1666464484
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1666464484
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1666464484
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1666464484
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1666464484
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1666464484
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1666464484
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1666464484
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1666464484
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1666464484
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1666464484
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1666464484
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1666464484
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1666464484
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1666464484
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1666464484
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1666464484
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1666464484
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1666464484
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1666464484
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1666464484
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1666464484
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1666464484
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1666464484
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_293
timestamp 1666464484
transform 1 0 28060 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_297
timestamp 1666464484
transform 1 0 28428 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1666464484
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_8
timestamp 1666464484
transform 1 0 1840 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_20
timestamp 1666464484
transform 1 0 2944 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1666464484
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1666464484
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1666464484
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1666464484
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1666464484
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1666464484
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1666464484
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1666464484
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1666464484
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1666464484
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1666464484
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1666464484
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1666464484
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1666464484
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1666464484
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1666464484
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1666464484
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1666464484
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1666464484
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1666464484
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1666464484
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1666464484
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1666464484
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1666464484
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1666464484
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1666464484
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1666464484
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_289
timestamp 1666464484
transform 1 0 27692 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_293
timestamp 1666464484
transform 1 0 28060 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_297
timestamp 1666464484
transform 1 0 28428 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1666464484
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_8
timestamp 1666464484
transform 1 0 1840 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_20
timestamp 1666464484
transform 1 0 2944 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_32
timestamp 1666464484
transform 1 0 4048 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_44
timestamp 1666464484
transform 1 0 5152 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1666464484
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1666464484
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1666464484
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1666464484
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1666464484
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1666464484
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1666464484
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1666464484
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1666464484
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1666464484
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1666464484
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1666464484
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1666464484
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1666464484
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1666464484
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1666464484
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1666464484
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1666464484
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1666464484
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1666464484
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1666464484
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1666464484
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1666464484
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1666464484
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1666464484
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_293
timestamp 1666464484
transform 1 0 28060 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1666464484
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1666464484
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1666464484
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1666464484
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1666464484
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1666464484
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1666464484
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1666464484
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1666464484
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1666464484
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1666464484
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1666464484
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1666464484
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1666464484
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1666464484
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1666464484
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1666464484
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1666464484
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1666464484
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1666464484
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1666464484
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1666464484
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1666464484
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1666464484
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1666464484
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1666464484
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1666464484
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1666464484
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1666464484
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1666464484
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_289
timestamp 1666464484
transform 1 0 27692 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_297
timestamp 1666464484
transform 1 0 28428 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1666464484
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1666464484
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1666464484
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1666464484
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1666464484
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1666464484
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1666464484
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1666464484
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1666464484
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1666464484
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1666464484
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1666464484
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1666464484
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1666464484
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1666464484
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1666464484
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1666464484
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1666464484
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1666464484
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1666464484
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1666464484
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1666464484
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1666464484
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1666464484
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1666464484
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1666464484
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1666464484
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1666464484
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1666464484
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1666464484
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1666464484
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_293
timestamp 1666464484
transform 1 0 28060 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_297
timestamp 1666464484
transform 1 0 28428 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1666464484
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_8
timestamp 1666464484
transform 1 0 1840 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_20
timestamp 1666464484
transform 1 0 2944 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1666464484
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1666464484
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1666464484
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1666464484
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1666464484
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1666464484
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1666464484
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1666464484
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1666464484
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1666464484
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1666464484
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1666464484
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1666464484
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1666464484
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1666464484
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1666464484
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1666464484
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1666464484
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1666464484
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1666464484
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1666464484
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1666464484
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1666464484
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1666464484
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1666464484
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1666464484
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1666464484
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_289
timestamp 1666464484
transform 1 0 27692 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_293
timestamp 1666464484
transform 1 0 28060 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_297
timestamp 1666464484
transform 1 0 28428 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1666464484
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_8
timestamp 1666464484
transform 1 0 1840 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_20
timestamp 1666464484
transform 1 0 2944 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_32
timestamp 1666464484
transform 1 0 4048 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_44
timestamp 1666464484
transform 1 0 5152 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1666464484
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1666464484
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1666464484
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1666464484
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1666464484
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1666464484
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1666464484
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1666464484
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1666464484
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1666464484
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1666464484
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1666464484
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1666464484
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1666464484
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1666464484
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1666464484
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1666464484
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1666464484
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1666464484
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1666464484
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1666464484
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1666464484
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1666464484
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1666464484
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1666464484
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_293
timestamp 1666464484
transform 1 0 28060 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1666464484
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1666464484
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1666464484
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1666464484
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1666464484
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1666464484
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1666464484
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1666464484
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1666464484
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1666464484
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1666464484
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1666464484
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1666464484
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1666464484
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1666464484
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1666464484
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1666464484
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1666464484
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1666464484
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1666464484
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1666464484
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1666464484
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1666464484
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1666464484
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1666464484
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1666464484
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1666464484
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1666464484
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1666464484
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1666464484
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_289
timestamp 1666464484
transform 1 0 27692 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_297
timestamp 1666464484
transform 1 0 28428 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1666464484
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_8
timestamp 1666464484
transform 1 0 1840 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_20
timestamp 1666464484
transform 1 0 2944 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_32
timestamp 1666464484
transform 1 0 4048 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_44
timestamp 1666464484
transform 1 0 5152 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1666464484
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1666464484
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1666464484
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1666464484
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1666464484
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1666464484
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1666464484
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1666464484
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1666464484
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1666464484
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1666464484
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1666464484
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1666464484
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1666464484
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1666464484
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1666464484
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1666464484
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1666464484
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1666464484
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1666464484
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1666464484
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1666464484
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1666464484
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1666464484
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1666464484
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_293
timestamp 1666464484
transform 1 0 28060 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_297
timestamp 1666464484
transform 1 0 28428 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1666464484
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1666464484
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1666464484
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1666464484
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1666464484
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1666464484
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1666464484
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1666464484
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1666464484
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1666464484
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1666464484
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1666464484
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1666464484
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1666464484
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1666464484
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1666464484
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1666464484
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1666464484
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1666464484
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1666464484
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1666464484
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1666464484
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1666464484
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1666464484
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1666464484
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1666464484
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1666464484
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1666464484
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1666464484
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1666464484
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_289
timestamp 1666464484
transform 1 0 27692 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_293
timestamp 1666464484
transform 1 0 28060 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_297
timestamp 1666464484
transform 1 0 28428 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1666464484
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_8
timestamp 1666464484
transform 1 0 1840 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_20
timestamp 1666464484
transform 1 0 2944 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_32
timestamp 1666464484
transform 1 0 4048 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_44
timestamp 1666464484
transform 1 0 5152 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1666464484
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1666464484
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1666464484
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1666464484
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1666464484
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1666464484
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1666464484
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1666464484
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1666464484
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1666464484
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1666464484
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1666464484
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1666464484
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1666464484
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1666464484
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1666464484
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1666464484
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1666464484
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1666464484
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1666464484
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1666464484
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1666464484
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1666464484
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1666464484
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1666464484
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_293
timestamp 1666464484
transform 1 0 28060 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1666464484
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1666464484
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1666464484
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1666464484
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1666464484
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1666464484
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1666464484
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1666464484
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1666464484
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_85
timestamp 1666464484
transform 1 0 8924 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_93
timestamp 1666464484
transform 1 0 9660 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_105
timestamp 1666464484
transform 1 0 10764 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_117
timestamp 1666464484
transform 1 0 11868 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_129
timestamp 1666464484
transform 1 0 12972 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_137
timestamp 1666464484
transform 1 0 13708 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1666464484
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1666464484
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1666464484
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1666464484
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1666464484
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1666464484
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1666464484
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1666464484
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1666464484
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1666464484
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1666464484
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1666464484
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1666464484
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1666464484
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1666464484
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_289
timestamp 1666464484
transform 1 0 27692 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_293
timestamp 1666464484
transform 1 0 28060 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_297
timestamp 1666464484
transform 1 0 28428 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1666464484
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_8
timestamp 1666464484
transform 1 0 1840 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_20
timestamp 1666464484
transform 1 0 2944 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_32
timestamp 1666464484
transform 1 0 4048 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_36
timestamp 1666464484
transform 1 0 4416 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_48
timestamp 1666464484
transform 1 0 5520 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_57
timestamp 1666464484
transform 1 0 6348 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_61
timestamp 1666464484
transform 1 0 6716 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_64
timestamp 1666464484
transform 1 0 6992 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_76
timestamp 1666464484
transform 1 0 8096 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_84
timestamp 1666464484
transform 1 0 8832 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_90
timestamp 1666464484
transform 1 0 9384 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_97
timestamp 1666464484
transform 1 0 10028 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_103
timestamp 1666464484
transform 1 0 10580 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_109
timestamp 1666464484
transform 1 0 11132 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1666464484
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1666464484
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1666464484
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1666464484
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1666464484
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1666464484
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1666464484
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1666464484
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1666464484
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1666464484
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1666464484
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1666464484
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1666464484
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1666464484
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1666464484
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1666464484
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1666464484
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1666464484
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1666464484
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_293
timestamp 1666464484
transform 1 0 28060 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1666464484
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_8
timestamp 1666464484
transform 1 0 1840 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_16
timestamp 1666464484
transform 1 0 2576 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_29
timestamp 1666464484
transform 1 0 3772 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_33
timestamp 1666464484
transform 1 0 4140 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_36
timestamp 1666464484
transform 1 0 4416 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_44
timestamp 1666464484
transform 1 0 5152 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_56
timestamp 1666464484
transform 1 0 6256 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_59
timestamp 1666464484
transform 1 0 6532 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_63
timestamp 1666464484
transform 1 0 6900 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_66
timestamp 1666464484
transform 1 0 7176 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_74
timestamp 1666464484
transform 1 0 7912 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_78
timestamp 1666464484
transform 1 0 8280 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1666464484
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1666464484
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_91
timestamp 1666464484
transform 1 0 9476 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_99
timestamp 1666464484
transform 1 0 10212 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_106
timestamp 1666464484
transform 1 0 10856 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_112
timestamp 1666464484
transform 1 0 11408 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_122
timestamp 1666464484
transform 1 0 12328 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_134
timestamp 1666464484
transform 1 0 13432 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1666464484
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1666464484
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1666464484
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1666464484
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1666464484
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1666464484
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1666464484
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1666464484
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1666464484
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1666464484
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1666464484
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1666464484
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1666464484
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1666464484
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1666464484
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_289
timestamp 1666464484
transform 1 0 27692 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_293
timestamp 1666464484
transform 1 0 28060 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_297
timestamp 1666464484
transform 1 0 28428 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_3
timestamp 1666464484
transform 1 0 1380 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_9
timestamp 1666464484
transform 1 0 1932 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_12
timestamp 1666464484
transform 1 0 2208 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_18
timestamp 1666464484
transform 1 0 2760 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_26
timestamp 1666464484
transform 1 0 3496 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_32
timestamp 1666464484
transform 1 0 4048 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_38
timestamp 1666464484
transform 1 0 4600 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_41_46
timestamp 1666464484
transform 1 0 5336 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_54
timestamp 1666464484
transform 1 0 6072 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_57
timestamp 1666464484
transform 1 0 6348 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_64
timestamp 1666464484
transform 1 0 6992 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_68
timestamp 1666464484
transform 1 0 7360 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_73
timestamp 1666464484
transform 1 0 7820 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_82
timestamp 1666464484
transform 1 0 8648 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_93
timestamp 1666464484
transform 1 0 9660 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_99
timestamp 1666464484
transform 1 0 10212 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_107
timestamp 1666464484
transform 1 0 10948 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1666464484
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 1666464484
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_119
timestamp 1666464484
transform 1 0 12052 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_125
timestamp 1666464484
transform 1 0 12604 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_131
timestamp 1666464484
transform 1 0 13156 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_134
timestamp 1666464484
transform 1 0 13432 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_146
timestamp 1666464484
transform 1 0 14536 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_158
timestamp 1666464484
transform 1 0 15640 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1666464484
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1666464484
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1666464484
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1666464484
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1666464484
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1666464484
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1666464484
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1666464484
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1666464484
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1666464484
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1666464484
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1666464484
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1666464484
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1666464484
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_293
timestamp 1666464484
transform 1 0 28060 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1666464484
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_8
timestamp 1666464484
transform 1 0 1840 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_15
timestamp 1666464484
transform 1 0 2484 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_23
timestamp 1666464484
transform 1 0 3220 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_26
timestamp 1666464484
transform 1 0 3496 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_29
timestamp 1666464484
transform 1 0 3772 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_33
timestamp 1666464484
transform 1 0 4140 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_36
timestamp 1666464484
transform 1 0 4416 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_42
timestamp 1666464484
transform 1 0 4968 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_46
timestamp 1666464484
transform 1 0 5336 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_49
timestamp 1666464484
transform 1 0 5612 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_56
timestamp 1666464484
transform 1 0 6256 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_64
timestamp 1666464484
transform 1 0 6992 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_72
timestamp 1666464484
transform 1 0 7728 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_82
timestamp 1666464484
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_85
timestamp 1666464484
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_89
timestamp 1666464484
transform 1 0 9292 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_93
timestamp 1666464484
transform 1 0 9660 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_99
timestamp 1666464484
transform 1 0 10212 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_108
timestamp 1666464484
transform 1 0 11040 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_114
timestamp 1666464484
transform 1 0 11592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_120
timestamp 1666464484
transform 1 0 12144 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_128
timestamp 1666464484
transform 1 0 12880 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_134
timestamp 1666464484
transform 1 0 13432 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1666464484
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_145
timestamp 1666464484
transform 1 0 14444 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_157
timestamp 1666464484
transform 1 0 15548 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_169
timestamp 1666464484
transform 1 0 16652 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_181
timestamp 1666464484
transform 1 0 17756 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_193
timestamp 1666464484
transform 1 0 18860 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1666464484
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1666464484
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1666464484
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1666464484
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1666464484
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1666464484
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1666464484
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1666464484
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1666464484
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_289
timestamp 1666464484
transform 1 0 27692 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_293
timestamp 1666464484
transform 1 0 28060 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_297
timestamp 1666464484
transform 1 0 28428 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_3
timestamp 1666464484
transform 1 0 1380 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_9
timestamp 1666464484
transform 1 0 1932 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_16
timestamp 1666464484
transform 1 0 2576 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_23
timestamp 1666464484
transform 1 0 3220 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_43_34
timestamp 1666464484
transform 1 0 4232 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_40
timestamp 1666464484
transform 1 0 4784 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_44
timestamp 1666464484
transform 1 0 5152 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_43_54
timestamp 1666464484
transform 1 0 6072 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_57
timestamp 1666464484
transform 1 0 6348 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_61
timestamp 1666464484
transform 1 0 6716 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_69
timestamp 1666464484
transform 1 0 7452 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_93
timestamp 1666464484
transform 1 0 9660 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_103
timestamp 1666464484
transform 1 0 10580 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_109
timestamp 1666464484
transform 1 0 11132 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_113
timestamp 1666464484
transform 1 0 11500 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_121
timestamp 1666464484
transform 1 0 12236 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_130
timestamp 1666464484
transform 1 0 13064 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_137
timestamp 1666464484
transform 1 0 13708 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_143
timestamp 1666464484
transform 1 0 14260 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1666464484
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1666464484
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1666464484
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_169
timestamp 1666464484
transform 1 0 16652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_175
timestamp 1666464484
transform 1 0 17204 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1666464484
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1666464484
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1666464484
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1666464484
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1666464484
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1666464484
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1666464484
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1666464484
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1666464484
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1666464484
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1666464484
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1666464484
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_293
timestamp 1666464484
transform 1 0 28060 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_297
timestamp 1666464484
transform 1 0 28428 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1666464484
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_8
timestamp 1666464484
transform 1 0 1840 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_16
timestamp 1666464484
transform 1 0 2576 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_24
timestamp 1666464484
transform 1 0 3312 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_29
timestamp 1666464484
transform 1 0 3772 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_34
timestamp 1666464484
transform 1 0 4232 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_42
timestamp 1666464484
transform 1 0 4968 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_54
timestamp 1666464484
transform 1 0 6072 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_62
timestamp 1666464484
transform 1 0 6808 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_74
timestamp 1666464484
transform 1 0 7912 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_82
timestamp 1666464484
transform 1 0 8648 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1666464484
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_103
timestamp 1666464484
transform 1 0 10580 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_111
timestamp 1666464484
transform 1 0 11316 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_121
timestamp 1666464484
transform 1 0 12236 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_130
timestamp 1666464484
transform 1 0 13064 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_138
timestamp 1666464484
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_141
timestamp 1666464484
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_146
timestamp 1666464484
transform 1 0 14536 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_152
timestamp 1666464484
transform 1 0 15088 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_158
timestamp 1666464484
transform 1 0 15640 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_170
timestamp 1666464484
transform 1 0 16744 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_182
timestamp 1666464484
transform 1 0 17848 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_194
timestamp 1666464484
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1666464484
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1666464484
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1666464484
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1666464484
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1666464484
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1666464484
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1666464484
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1666464484
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1666464484
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_289
timestamp 1666464484
transform 1 0 27692 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_297
timestamp 1666464484
transform 1 0 28428 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1666464484
transform 1 0 1380 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_9
timestamp 1666464484
transform 1 0 1932 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_17
timestamp 1666464484
transform 1 0 2668 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_21
timestamp 1666464484
transform 1 0 3036 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_26
timestamp 1666464484
transform 1 0 3496 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_33
timestamp 1666464484
transform 1 0 4140 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_37
timestamp 1666464484
transform 1 0 4508 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_54
timestamp 1666464484
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_57
timestamp 1666464484
transform 1 0 6348 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_75
timestamp 1666464484
transform 1 0 8004 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_84
timestamp 1666464484
transform 1 0 8832 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_104
timestamp 1666464484
transform 1 0 10672 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_110
timestamp 1666464484
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_113
timestamp 1666464484
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_125
timestamp 1666464484
transform 1 0 12604 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_135
timestamp 1666464484
transform 1 0 13524 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_144
timestamp 1666464484
transform 1 0 14352 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_152
timestamp 1666464484
transform 1 0 15088 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_160
timestamp 1666464484
transform 1 0 15824 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 1666464484
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1666464484
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1666464484
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1666464484
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1666464484
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1666464484
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1666464484
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1666464484
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1666464484
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1666464484
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1666464484
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1666464484
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1666464484
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1666464484
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_293
timestamp 1666464484
transform 1 0 28060 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_46_3
timestamp 1666464484
transform 1 0 1380 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_14
timestamp 1666464484
transform 1 0 2392 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_26
timestamp 1666464484
transform 1 0 3496 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_29
timestamp 1666464484
transform 1 0 3772 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_41
timestamp 1666464484
transform 1 0 4876 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_45
timestamp 1666464484
transform 1 0 5244 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_62
timestamp 1666464484
transform 1 0 6808 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_82
timestamp 1666464484
transform 1 0 8648 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_85
timestamp 1666464484
transform 1 0 8924 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_105
timestamp 1666464484
transform 1 0 10764 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_111
timestamp 1666464484
transform 1 0 11316 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_125
timestamp 1666464484
transform 1 0 12604 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_135
timestamp 1666464484
transform 1 0 13524 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1666464484
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_141
timestamp 1666464484
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_148
timestamp 1666464484
transform 1 0 14720 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_157
timestamp 1666464484
transform 1 0 15548 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_165
timestamp 1666464484
transform 1 0 16284 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_172
timestamp 1666464484
transform 1 0 16928 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_178
timestamp 1666464484
transform 1 0 17480 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_190
timestamp 1666464484
transform 1 0 18584 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1666464484
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1666464484
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1666464484
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1666464484
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1666464484
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1666464484
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1666464484
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1666464484
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1666464484
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_289
timestamp 1666464484
transform 1 0 27692 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_293
timestamp 1666464484
transform 1 0 28060 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_297
timestamp 1666464484
transform 1 0 28428 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_3
timestamp 1666464484
transform 1 0 1380 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_9
timestamp 1666464484
transform 1 0 1932 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_26
timestamp 1666464484
transform 1 0 3496 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_34
timestamp 1666464484
transform 1 0 4232 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_54
timestamp 1666464484
transform 1 0 6072 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_57
timestamp 1666464484
transform 1 0 6348 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_66
timestamp 1666464484
transform 1 0 7176 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_86
timestamp 1666464484
transform 1 0 9016 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_106
timestamp 1666464484
transform 1 0 10856 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_113
timestamp 1666464484
transform 1 0 11500 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_131
timestamp 1666464484
transform 1 0 13156 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_145
timestamp 1666464484
transform 1 0 14444 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_155
timestamp 1666464484
transform 1 0 15364 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_164
timestamp 1666464484
transform 1 0 16192 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_169
timestamp 1666464484
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_173
timestamp 1666464484
transform 1 0 17020 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_185
timestamp 1666464484
transform 1 0 18124 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_197
timestamp 1666464484
transform 1 0 19228 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_209
timestamp 1666464484
transform 1 0 20332 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_221
timestamp 1666464484
transform 1 0 21436 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1666464484
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1666464484
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1666464484
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1666464484
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1666464484
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1666464484
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1666464484
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_293
timestamp 1666464484
transform 1 0 28060 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_297
timestamp 1666464484
transform 1 0 28428 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_3
timestamp 1666464484
transform 1 0 1380 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_9
timestamp 1666464484
transform 1 0 1932 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_26
timestamp 1666464484
transform 1 0 3496 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_29
timestamp 1666464484
transform 1 0 3772 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_41
timestamp 1666464484
transform 1 0 4876 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_65
timestamp 1666464484
transform 1 0 7084 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_76
timestamp 1666464484
transform 1 0 8096 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_82
timestamp 1666464484
transform 1 0 8648 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_85
timestamp 1666464484
transform 1 0 8924 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_97
timestamp 1666464484
transform 1 0 10028 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_105
timestamp 1666464484
transform 1 0 10764 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_126
timestamp 1666464484
transform 1 0 12696 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_48_137
timestamp 1666464484
transform 1 0 13708 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_141
timestamp 1666464484
transform 1 0 14076 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_151
timestamp 1666464484
transform 1 0 14996 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_161
timestamp 1666464484
transform 1 0 15916 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_169
timestamp 1666464484
transform 1 0 16652 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_176
timestamp 1666464484
transform 1 0 17296 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_182
timestamp 1666464484
transform 1 0 17848 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_188
timestamp 1666464484
transform 1 0 18400 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1666464484
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1666464484
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1666464484
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1666464484
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1666464484
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1666464484
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1666464484
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1666464484
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1666464484
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_289
timestamp 1666464484
transform 1 0 27692 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_297
timestamp 1666464484
transform 1 0 28428 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_3
timestamp 1666464484
transform 1 0 1380 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_7
timestamp 1666464484
transform 1 0 1748 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_14
timestamp 1666464484
transform 1 0 2392 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_34
timestamp 1666464484
transform 1 0 4232 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_54
timestamp 1666464484
transform 1 0 6072 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_57
timestamp 1666464484
transform 1 0 6348 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_69
timestamp 1666464484
transform 1 0 7452 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_93
timestamp 1666464484
transform 1 0 9660 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_99
timestamp 1666464484
transform 1 0 10212 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_107
timestamp 1666464484
transform 1 0 10948 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_110
timestamp 1666464484
transform 1 0 11224 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_113
timestamp 1666464484
transform 1 0 11500 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_117
timestamp 1666464484
transform 1 0 11868 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_125
timestamp 1666464484
transform 1 0 12604 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_149
timestamp 1666464484
transform 1 0 14812 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_163
timestamp 1666464484
transform 1 0 16100 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1666464484
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1666464484
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_175
timestamp 1666464484
transform 1 0 17204 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_182
timestamp 1666464484
transform 1 0 17848 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_188
timestamp 1666464484
transform 1 0 18400 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_200
timestamp 1666464484
transform 1 0 19504 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_212
timestamp 1666464484
transform 1 0 20608 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1666464484
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1666464484
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1666464484
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1666464484
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1666464484
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1666464484
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1666464484
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_293
timestamp 1666464484
transform 1 0 28060 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_50_3
timestamp 1666464484
transform 1 0 1380 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_9
timestamp 1666464484
transform 1 0 1932 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_26
timestamp 1666464484
transform 1 0 3496 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_29
timestamp 1666464484
transform 1 0 3772 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_42
timestamp 1666464484
transform 1 0 4968 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_62
timestamp 1666464484
transform 1 0 6808 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_82
timestamp 1666464484
transform 1 0 8648 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_85
timestamp 1666464484
transform 1 0 8924 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_89
timestamp 1666464484
transform 1 0 9292 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_106
timestamp 1666464484
transform 1 0 10856 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_114
timestamp 1666464484
transform 1 0 11592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_131
timestamp 1666464484
transform 1 0 13156 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_135
timestamp 1666464484
transform 1 0 13524 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_138
timestamp 1666464484
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_141
timestamp 1666464484
transform 1 0 14076 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_150
timestamp 1666464484
transform 1 0 14904 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_160
timestamp 1666464484
transform 1 0 15824 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_170
timestamp 1666464484
transform 1 0 16744 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_179
timestamp 1666464484
transform 1 0 17572 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_187
timestamp 1666464484
transform 1 0 18308 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_194
timestamp 1666464484
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_197
timestamp 1666464484
transform 1 0 19228 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_201
timestamp 1666464484
transform 1 0 19596 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_207
timestamp 1666464484
transform 1 0 20148 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_213
timestamp 1666464484
transform 1 0 20700 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_225
timestamp 1666464484
transform 1 0 21804 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_237
timestamp 1666464484
transform 1 0 22908 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_249
timestamp 1666464484
transform 1 0 24012 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1666464484
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1666464484
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1666464484
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_289
timestamp 1666464484
transform 1 0 27692 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_293
timestamp 1666464484
transform 1 0 28060 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_297
timestamp 1666464484
transform 1 0 28428 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_3
timestamp 1666464484
transform 1 0 1380 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_7
timestamp 1666464484
transform 1 0 1748 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_14
timestamp 1666464484
transform 1 0 2392 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_34
timestamp 1666464484
transform 1 0 4232 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_54
timestamp 1666464484
transform 1 0 6072 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_57
timestamp 1666464484
transform 1 0 6348 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_63
timestamp 1666464484
transform 1 0 6900 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_87
timestamp 1666464484
transform 1 0 9108 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_107
timestamp 1666464484
transform 1 0 10948 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1666464484
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_113
timestamp 1666464484
transform 1 0 11500 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_131
timestamp 1666464484
transform 1 0 13156 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_151
timestamp 1666464484
transform 1 0 14996 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_162
timestamp 1666464484
transform 1 0 16008 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_51_169
timestamp 1666464484
transform 1 0 16652 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_177
timestamp 1666464484
transform 1 0 17388 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_186
timestamp 1666464484
transform 1 0 18216 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_194
timestamp 1666464484
transform 1 0 18952 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_201
timestamp 1666464484
transform 1 0 19596 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_207
timestamp 1666464484
transform 1 0 20148 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_213
timestamp 1666464484
transform 1 0 20700 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_221
timestamp 1666464484
transform 1 0 21436 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1666464484
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1666464484
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1666464484
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1666464484
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1666464484
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1666464484
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1666464484
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_293
timestamp 1666464484
transform 1 0 28060 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_297
timestamp 1666464484
transform 1 0 28428 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_3
timestamp 1666464484
transform 1 0 1380 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_9
timestamp 1666464484
transform 1 0 1932 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_26
timestamp 1666464484
transform 1 0 3496 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_29
timestamp 1666464484
transform 1 0 3772 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_42
timestamp 1666464484
transform 1 0 4968 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_62
timestamp 1666464484
transform 1 0 6808 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_82
timestamp 1666464484
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_85
timestamp 1666464484
transform 1 0 8924 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_90
timestamp 1666464484
transform 1 0 9384 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_110
timestamp 1666464484
transform 1 0 11224 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_117
timestamp 1666464484
transform 1 0 11868 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_52_137
timestamp 1666464484
transform 1 0 13708 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_141
timestamp 1666464484
transform 1 0 14076 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_159
timestamp 1666464484
transform 1 0 15732 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_170
timestamp 1666464484
transform 1 0 16744 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_180
timestamp 1666464484
transform 1 0 17664 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1666464484
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1666464484
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_197
timestamp 1666464484
transform 1 0 19228 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_203
timestamp 1666464484
transform 1 0 19780 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_210
timestamp 1666464484
transform 1 0 20424 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_216
timestamp 1666464484
transform 1 0 20976 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_222
timestamp 1666464484
transform 1 0 21528 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_234
timestamp 1666464484
transform 1 0 22632 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_246
timestamp 1666464484
transform 1 0 23736 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1666464484
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1666464484
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_277
timestamp 1666464484
transform 1 0 26588 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_285
timestamp 1666464484
transform 1 0 27324 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_290
timestamp 1666464484
transform 1 0 27784 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_297
timestamp 1666464484
transform 1 0 28428 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_3
timestamp 1666464484
transform 1 0 1380 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_9
timestamp 1666464484
transform 1 0 1932 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_26
timestamp 1666464484
transform 1 0 3496 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_29
timestamp 1666464484
transform 1 0 3772 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_34
timestamp 1666464484
transform 1 0 4232 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_54
timestamp 1666464484
transform 1 0 6072 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_57
timestamp 1666464484
transform 1 0 6348 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_62
timestamp 1666464484
transform 1 0 6808 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_82
timestamp 1666464484
transform 1 0 8648 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_85
timestamp 1666464484
transform 1 0 8924 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_90
timestamp 1666464484
transform 1 0 9384 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_110
timestamp 1666464484
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_113
timestamp 1666464484
transform 1 0 11500 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_131
timestamp 1666464484
transform 1 0 13156 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_137
timestamp 1666464484
transform 1 0 13708 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_141
timestamp 1666464484
transform 1 0 14076 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_159
timestamp 1666464484
transform 1 0 15732 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_166
timestamp 1666464484
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_169
timestamp 1666464484
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_187
timestamp 1666464484
transform 1 0 18308 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_194
timestamp 1666464484
transform 1 0 18952 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_197
timestamp 1666464484
transform 1 0 19228 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_204
timestamp 1666464484
transform 1 0 19872 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_212
timestamp 1666464484
transform 1 0 20608 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_219
timestamp 1666464484
transform 1 0 21252 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1666464484
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_225
timestamp 1666464484
transform 1 0 21804 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_230
timestamp 1666464484
transform 1 0 22264 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_242
timestamp 1666464484
transform 1 0 23368 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_246
timestamp 1666464484
transform 1 0 23736 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_250
timestamp 1666464484
transform 1 0 24104 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_253
timestamp 1666464484
transform 1 0 24380 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_262
timestamp 1666464484
transform 1 0 25208 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_274
timestamp 1666464484
transform 1 0 26312 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_281
timestamp 1666464484
transform 1 0 26956 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_286
timestamp 1666464484
transform 1 0 27416 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_297
timestamp 1666464484
transform 1 0 28428 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666464484
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666464484
transform -1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666464484
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666464484
transform -1 0 28888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666464484
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666464484
transform -1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666464484
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666464484
transform -1 0 28888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666464484
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666464484
transform -1 0 28888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666464484
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666464484
transform -1 0 28888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666464484
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666464484
transform -1 0 28888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666464484
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666464484
transform -1 0 28888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666464484
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666464484
transform -1 0 28888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666464484
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666464484
transform -1 0 28888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666464484
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666464484
transform -1 0 28888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666464484
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666464484
transform -1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666464484
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666464484
transform -1 0 28888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666464484
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666464484
transform -1 0 28888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666464484
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666464484
transform -1 0 28888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666464484
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666464484
transform -1 0 28888 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666464484
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666464484
transform -1 0 28888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666464484
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666464484
transform -1 0 28888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666464484
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666464484
transform -1 0 28888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666464484
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666464484
transform -1 0 28888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666464484
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666464484
transform -1 0 28888 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666464484
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666464484
transform -1 0 28888 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666464484
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666464484
transform -1 0 28888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666464484
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666464484
transform -1 0 28888 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666464484
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666464484
transform -1 0 28888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1666464484
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1666464484
transform -1 0 28888 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1666464484
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1666464484
transform -1 0 28888 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1666464484
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1666464484
transform -1 0 28888 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1666464484
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1666464484
transform -1 0 28888 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1666464484
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1666464484
transform -1 0 28888 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1666464484
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1666464484
transform -1 0 28888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1666464484
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1666464484
transform -1 0 28888 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1666464484
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1666464484
transform -1 0 28888 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1666464484
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1666464484
transform -1 0 28888 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1666464484
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1666464484
transform -1 0 28888 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1666464484
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1666464484
transform -1 0 28888 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1666464484
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1666464484
transform -1 0 28888 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1666464484
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1666464484
transform -1 0 28888 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1666464484
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1666464484
transform -1 0 28888 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1666464484
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1666464484
transform -1 0 28888 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1666464484
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1666464484
transform -1 0 28888 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1666464484
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1666464484
transform -1 0 28888 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1666464484
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1666464484
transform -1 0 28888 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1666464484
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1666464484
transform -1 0 28888 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1666464484
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1666464484
transform -1 0 28888 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1666464484
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1666464484
transform -1 0 28888 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1666464484
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1666464484
transform -1 0 28888 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1666464484
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1666464484
transform -1 0 28888 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1666464484
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1666464484
transform -1 0 28888 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1666464484
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1666464484
transform -1 0 28888 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1666464484
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1666464484
transform -1 0 28888 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1666464484
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1666464484
transform -1 0 28888 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1666464484
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1666464484
transform -1 0 28888 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1666464484
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1666464484
transform -1 0 28888 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1666464484
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1666464484
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1666464484
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1666464484
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1666464484
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1666464484
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1666464484
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1666464484
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1666464484
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1666464484
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1666464484
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1666464484
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1666464484
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1666464484
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1666464484
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1666464484
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1666464484
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1666464484
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1666464484
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1666464484
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1666464484
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1666464484
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1666464484
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1666464484
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1666464484
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1666464484
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1666464484
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1666464484
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1666464484
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1666464484
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1666464484
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1666464484
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1666464484
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1666464484
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1666464484
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1666464484
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1666464484
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1666464484
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1666464484
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1666464484
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1666464484
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1666464484
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1666464484
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1666464484
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1666464484
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1666464484
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1666464484
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1666464484
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1666464484
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1666464484
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1666464484
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1666464484
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1666464484
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1666464484
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1666464484
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1666464484
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1666464484
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1666464484
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1666464484
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1666464484
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1666464484
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1666464484
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1666464484
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1666464484
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1666464484
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1666464484
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1666464484
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1666464484
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1666464484
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1666464484
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1666464484
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1666464484
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1666464484
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1666464484
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1666464484
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1666464484
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1666464484
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1666464484
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1666464484
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1666464484
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1666464484
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1666464484
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1666464484
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1666464484
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1666464484
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1666464484
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1666464484
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1666464484
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1666464484
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1666464484
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1666464484
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1666464484
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1666464484
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1666464484
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1666464484
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1666464484
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1666464484
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1666464484
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1666464484
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1666464484
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1666464484
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1666464484
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1666464484
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1666464484
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1666464484
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1666464484
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1666464484
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1666464484
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1666464484
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1666464484
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1666464484
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1666464484
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1666464484
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1666464484
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1666464484
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1666464484
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1666464484
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1666464484
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1666464484
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1666464484
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1666464484
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1666464484
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1666464484
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1666464484
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1666464484
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1666464484
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1666464484
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1666464484
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1666464484
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1666464484
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1666464484
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1666464484
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1666464484
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1666464484
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1666464484
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1666464484
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1666464484
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1666464484
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1666464484
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1666464484
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1666464484
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1666464484
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1666464484
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1666464484
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1666464484
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1666464484
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1666464484
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1666464484
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1666464484
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1666464484
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1666464484
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1666464484
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1666464484
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1666464484
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1666464484
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1666464484
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1666464484
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1666464484
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1666464484
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1666464484
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1666464484
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1666464484
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1666464484
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1666464484
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1666464484
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1666464484
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1666464484
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1666464484
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1666464484
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1666464484
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1666464484
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1666464484
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1666464484
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1666464484
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1666464484
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1666464484
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1666464484
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1666464484
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1666464484
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1666464484
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1666464484
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1666464484
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1666464484
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1666464484
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1666464484
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1666464484
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1666464484
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1666464484
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1666464484
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1666464484
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1666464484
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1666464484
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1666464484
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1666464484
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1666464484
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1666464484
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1666464484
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1666464484
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1666464484
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1666464484
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1666464484
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1666464484
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1666464484
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1666464484
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1666464484
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1666464484
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1666464484
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1666464484
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1666464484
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1666464484
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1666464484
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1666464484
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1666464484
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1666464484
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1666464484
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1666464484
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1666464484
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1666464484
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1666464484
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1666464484
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1666464484
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1666464484
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1666464484
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1666464484
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1666464484
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1666464484
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1666464484
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1666464484
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1666464484
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1666464484
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1666464484
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1666464484
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1666464484
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1666464484
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1666464484
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1666464484
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1666464484
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1666464484
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1666464484
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1666464484
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1666464484
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1666464484
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1666464484
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1666464484
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1666464484
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1666464484
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1666464484
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1666464484
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1666464484
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1666464484
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1666464484
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1666464484
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1666464484
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1666464484
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1666464484
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1666464484
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1666464484
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1666464484
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1666464484
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1666464484
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1666464484
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1666464484
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1666464484
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1666464484
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1666464484
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1666464484
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1666464484
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1666464484
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1666464484
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1666464484
transform 1 0 3680 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1666464484
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1666464484
transform 1 0 8832 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1666464484
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1666464484
transform 1 0 13984 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1666464484
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1666464484
transform 1 0 19136 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1666464484
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1666464484
transform 1 0 24288 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1666464484
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _093_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 17204 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _094_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 4232 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _095_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 14720 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _096_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5980 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _097_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 4232 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _098_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 16100 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _099_
timestamp 1666464484
transform -1 0 9384 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _100_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 20240 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _101_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 18492 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _102_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 13800 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _103_
timestamp 1666464484
transform 1 0 12512 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _104_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 14996 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _105_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 9384 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _106_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 15364 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _107_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 11684 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _108_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 10580 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _109_
timestamp 1666464484
transform -1 0 10856 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _110_
timestamp 1666464484
transform 1 0 19412 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _111_
timestamp 1666464484
transform 1 0 20148 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _112_
timestamp 1666464484
transform 1 0 16192 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _113_
timestamp 1666464484
transform -1 0 18216 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _114_
timestamp 1666464484
transform 1 0 17572 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _115_
timestamp 1666464484
transform 1 0 11684 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _116_
timestamp 1666464484
transform -1 0 11040 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _117_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 4968 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _118_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6532 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _119_
timestamp 1666464484
transform 1 0 8280 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _120_
timestamp 1666464484
transform 1 0 9752 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _121_
timestamp 1666464484
transform 1 0 15916 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _122_
timestamp 1666464484
transform 1 0 1840 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _123_
timestamp 1666464484
transform -1 0 3496 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _124_
timestamp 1666464484
transform 1 0 13892 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _125_
timestamp 1666464484
transform -1 0 6992 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _126_
timestamp 1666464484
transform -1 0 15088 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _127_
timestamp 1666464484
transform 1 0 13892 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _128_
timestamp 1666464484
transform 1 0 11684 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _129_
timestamp 1666464484
transform 1 0 8372 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _130_
timestamp 1666464484
transform -1 0 13708 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _131_
timestamp 1666464484
transform -1 0 3496 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _132_
timestamp 1666464484
transform 1 0 15732 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _133_
timestamp 1666464484
transform 1 0 16284 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _134_
timestamp 1666464484
transform 1 0 18676 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _135_
timestamp 1666464484
transform 1 0 12604 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _136_
timestamp 1666464484
transform 1 0 17020 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _137_
timestamp 1666464484
transform -1 0 10580 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _138_
timestamp 1666464484
transform -1 0 8096 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _139_
timestamp 1666464484
transform 1 0 19320 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _140_
timestamp 1666464484
transform -1 0 17388 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _141_
timestamp 1666464484
transform 1 0 9752 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _142_
timestamp 1666464484
transform 1 0 9844 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _143_
timestamp 1666464484
transform 1 0 16652 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _144_
timestamp 1666464484
transform -1 0 17572 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _145_
timestamp 1666464484
transform 1 0 14260 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _146_
timestamp 1666464484
transform 1 0 11684 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _147_
timestamp 1666464484
transform 1 0 15364 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _148_
timestamp 1666464484
transform -1 0 12604 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _149_
timestamp 1666464484
transform -1 0 4232 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _150_
timestamp 1666464484
transform 1 0 12972 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _151_
timestamp 1666464484
transform -1 0 6900 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _152_
timestamp 1666464484
transform 1 0 14812 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _153_
timestamp 1666464484
transform -1 0 7452 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _154_
timestamp 1666464484
transform -1 0 13064 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _155_
timestamp 1666464484
transform -1 0 3312 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _156_
timestamp 1666464484
transform -1 0 16744 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _157_
timestamp 1666464484
transform -1 0 12604 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _158_
timestamp 1666464484
transform -1 0 13708 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _159_
timestamp 1666464484
transform 1 0 17112 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _160_
timestamp 1666464484
transform -1 0 18308 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _161_
timestamp 1666464484
transform 1 0 15272 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _162_
timestamp 1666464484
transform 1 0 16836 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _163_
timestamp 1666464484
transform -1 0 15548 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _164_
timestamp 1666464484
transform 1 0 19412 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _165_
timestamp 1666464484
transform 1 0 14260 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _166_
timestamp 1666464484
transform -1 0 10028 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _167_
timestamp 1666464484
transform -1 0 6808 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _168_
timestamp 1666464484
transform 1 0 12972 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _169_
timestamp 1666464484
transform -1 0 2576 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _170_
timestamp 1666464484
transform 1 0 5520 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _171_
timestamp 1666464484
transform -1 0 6072 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _172_
timestamp 1666464484
transform -1 0 8648 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _173_
timestamp 1666464484
transform 1 0 1932 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _174_
timestamp 1666464484
transform 1 0 6440 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _175_
timestamp 1666464484
transform -1 0 9660 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _176_
timestamp 1666464484
transform 1 0 8372 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _177_
timestamp 1666464484
transform -1 0 8648 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _178_
timestamp 1666464484
transform -1 0 4968 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _179_
timestamp 1666464484
transform 1 0 6716 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _180_
timestamp 1666464484
transform 1 0 4324 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _181_
timestamp 1666464484
transform 1 0 7360 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _182_
timestamp 1666464484
transform -1 0 2392 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _183_
timestamp 1666464484
transform 1 0 9108 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _184_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6532 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _185_
timestamp 1666464484
transform -1 0 4140 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _186_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2760 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _187_
timestamp 1666464484
transform 1 0 4600 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _188_
timestamp 1666464484
transform -1 0 13156 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _189_
timestamp 1666464484
transform 1 0 14260 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _190_
timestamp 1666464484
transform 1 0 9752 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _191_
timestamp 1666464484
transform 1 0 7636 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _192_
timestamp 1666464484
transform 1 0 2024 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _193_
timestamp 1666464484
transform 1 0 2024 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _194_
timestamp 1666464484
transform -1 0 8004 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _195_
timestamp 1666464484
transform -1 0 6808 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _196_
timestamp 1666464484
transform -1 0 6072 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _197_
timestamp 1666464484
transform 1 0 9752 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _198_
timestamp 1666464484
transform 1 0 4600 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _199_
timestamp 1666464484
transform 1 0 11684 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _200_
timestamp 1666464484
transform -1 0 8648 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _201_
timestamp 1666464484
transform 1 0 2024 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _202_
timestamp 1666464484
transform -1 0 6808 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _203_
timestamp 1666464484
transform 1 0 2760 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _204_
timestamp 1666464484
transform 1 0 9200 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _205_
timestamp 1666464484
transform -1 0 10764 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _206_
timestamp 1666464484
transform 1 0 9384 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _207_
timestamp 1666464484
transform -1 0 6808 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _208_
timestamp 1666464484
transform -1 0 15732 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _209_
timestamp 1666464484
transform -1 0 14996 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _210_
timestamp 1666464484
transform -1 0 13156 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _211_
timestamp 1666464484
transform 1 0 4600 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _212_
timestamp 1666464484
transform 1 0 2024 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _213_
timestamp 1666464484
transform 1 0 11684 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _214_
timestamp 1666464484
transform 1 0 9476 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _215_
timestamp 1666464484
transform 1 0 9384 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _216_
timestamp 1666464484
transform 1 0 12236 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _217_
timestamp 1666464484
transform 1 0 7176 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _218_
timestamp 1666464484
transform 1 0 7176 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _219_
timestamp 1666464484
transform -1 0 3496 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _220_
timestamp 1666464484
transform 1 0 7544 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _221_
timestamp 1666464484
transform 1 0 9108 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _222_
timestamp 1666464484
transform 1 0 4600 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _223_
timestamp 1666464484
transform 1 0 16836 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _224_
timestamp 1666464484
transform 1 0 7176 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_io_in[0] pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 12696 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_io_in[0]
timestamp 1666464484
transform -1 0 9660 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_io_in[0]
timestamp 1666464484
transform -1 0 7084 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_io_in[0]
timestamp 1666464484
transform -1 0 9660 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_io_in[0]
timestamp 1666464484
transform 1 0 12972 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 7912 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1666464484
transform -1 0 4876 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1
timestamp 1666464484
transform -1 0 28428 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  output2
timestamp 1666464484
transform 1 0 18584 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp 1666464484
transform 1 0 12236 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 1666464484
transform 1 0 15456 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1666464484
transform 1 0 7452 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1666464484
transform 1 0 4600 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1666464484
transform -1 0 2668 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1666464484
transform -1 0 1932 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1666464484
transform -1 0 1932 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_10 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 1840 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_11
timestamp 1666464484
transform 1 0 28152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_12
timestamp 1666464484
transform 1 0 28152 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_13
timestamp 1666464484
transform 1 0 28152 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_14
timestamp 1666464484
transform 1 0 28152 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_15
timestamp 1666464484
transform 1 0 28152 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_16
timestamp 1666464484
transform 1 0 28152 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_17
timestamp 1666464484
transform 1 0 28152 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_18
timestamp 1666464484
transform 1 0 28152 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_19
timestamp 1666464484
transform 1 0 28152 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_20
timestamp 1666464484
transform 1 0 28152 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_21
timestamp 1666464484
transform 1 0 28152 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_22
timestamp 1666464484
transform 1 0 28152 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_23
timestamp 1666464484
transform 1 0 28152 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_24
timestamp 1666464484
transform 1 0 28152 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_25
timestamp 1666464484
transform 1 0 28152 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_26
timestamp 1666464484
transform -1 0 28428 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_27
timestamp 1666464484
transform -1 0 25208 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_28
timestamp 1666464484
transform -1 0 22264 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_29
timestamp 1666464484
transform -1 0 1840 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_30
timestamp 1666464484
transform -1 0 1840 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_31
timestamp 1666464484
transform -1 0 1840 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_32
timestamp 1666464484
transform -1 0 1840 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_33
timestamp 1666464484
transform -1 0 1840 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_34
timestamp 1666464484
transform -1 0 1840 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_35
timestamp 1666464484
transform -1 0 1840 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_36
timestamp 1666464484
transform -1 0 1840 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_37
timestamp 1666464484
transform -1 0 1840 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_38
timestamp 1666464484
transform -1 0 1840 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_39
timestamp 1666464484
transform -1 0 1840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_40
timestamp 1666464484
transform -1 0 1840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_41
timestamp 1666464484
transform 1 0 28152 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_42
timestamp 1666464484
transform 1 0 28152 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_43
timestamp 1666464484
transform 1 0 28152 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_44
timestamp 1666464484
transform 1 0 28152 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_45
timestamp 1666464484
transform 1 0 28152 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_46
timestamp 1666464484
transform 1 0 28152 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_47
timestamp 1666464484
transform 1 0 28152 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_48
timestamp 1666464484
transform 1 0 28152 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_49
timestamp 1666464484
transform 1 0 28152 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_50
timestamp 1666464484
transform 1 0 28152 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_51
timestamp 1666464484
transform 1 0 28152 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_52
timestamp 1666464484
transform 1 0 28152 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_53
timestamp 1666464484
transform 1 0 28152 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_54
timestamp 1666464484
transform 1 0 28152 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_55
timestamp 1666464484
transform 1 0 27508 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_56
timestamp 1666464484
transform -1 0 27416 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_57
timestamp 1666464484
transform -1 0 24104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_58
timestamp 1666464484
transform -1 0 21252 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_59
timestamp 1666464484
transform -1 0 18952 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_60
timestamp 1666464484
transform -1 0 16376 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_61
timestamp 1666464484
transform -1 0 11868 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_62
timestamp 1666464484
transform 1 0 4876 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_63
timestamp 1666464484
transform -1 0 4232 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_64
timestamp 1666464484
transform -1 0 3220 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_65
timestamp 1666464484
transform -1 0 2484 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_66
timestamp 1666464484
transform -1 0 1840 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_67
timestamp 1666464484
transform -1 0 2576 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_68
timestamp 1666464484
transform -1 0 1840 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_69
timestamp 1666464484
transform -1 0 1840 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_70
timestamp 1666464484
transform -1 0 1840 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_71
timestamp 1666464484
transform -1 0 1840 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_72
timestamp 1666464484
transform -1 0 1840 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_73
timestamp 1666464484
transform -1 0 1840 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_74
timestamp 1666464484
transform -1 0 1840 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_75
timestamp 1666464484
transform -1 0 1840 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_76
timestamp 1666464484
transform -1 0 1840 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_77
timestamp 1666464484
transform -1 0 1840 0 -1 5440
box -38 -48 314 592
<< labels >>
flabel metal3 s 29200 1912 30000 2032 0 FreeSans 480 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 29200 22312 30000 22432 0 FreeSans 480 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 29200 24352 30000 24472 0 FreeSans 480 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal3 s 29200 26392 30000 26512 0 FreeSans 480 0 0 0 io_in[12]
port 3 nsew signal input
flabel metal3 s 29200 28432 30000 28552 0 FreeSans 480 0 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 29200 30472 30000 30592 0 FreeSans 480 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 29274 33200 29330 34000 0 FreeSans 224 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 25962 33200 26018 34000 0 FreeSans 224 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 22650 33200 22706 34000 0 FreeSans 224 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 19338 33200 19394 34000 0 FreeSans 224 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 16026 33200 16082 34000 0 FreeSans 224 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 29200 3952 30000 4072 0 FreeSans 480 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 12714 33200 12770 34000 0 FreeSans 224 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 9402 33200 9458 34000 0 FreeSans 224 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 6090 33200 6146 34000 0 FreeSans 224 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 2778 33200 2834 34000 0 FreeSans 224 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s 0 30880 800 31000 0 FreeSans 480 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal3 s 0 28840 800 28960 0 FreeSans 480 0 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s 0 26800 800 26920 0 FreeSans 480 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s 0 24760 800 24880 0 FreeSans 480 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s 0 22720 800 22840 0 FreeSans 480 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s 0 20680 800 20800 0 FreeSans 480 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 29200 5992 30000 6112 0 FreeSans 480 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 io_in[31]
port 24 nsew signal input
flabel metal3 s 0 14560 800 14680 0 FreeSans 480 0 0 0 io_in[32]
port 25 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 io_in[33]
port 26 nsew signal input
flabel metal3 s 0 10480 800 10600 0 FreeSans 480 0 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 29200 8032 30000 8152 0 FreeSans 480 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal3 s 29200 10072 30000 10192 0 FreeSans 480 0 0 0 io_in[4]
port 32 nsew signal input
flabel metal3 s 29200 12112 30000 12232 0 FreeSans 480 0 0 0 io_in[5]
port 33 nsew signal input
flabel metal3 s 29200 14152 30000 14272 0 FreeSans 480 0 0 0 io_in[6]
port 34 nsew signal input
flabel metal3 s 29200 16192 30000 16312 0 FreeSans 480 0 0 0 io_in[7]
port 35 nsew signal input
flabel metal3 s 29200 18232 30000 18352 0 FreeSans 480 0 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 29200 20272 30000 20392 0 FreeSans 480 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal3 s 29200 3272 30000 3392 0 FreeSans 480 0 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 29200 23672 30000 23792 0 FreeSans 480 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 29200 25712 30000 25832 0 FreeSans 480 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal3 s 29200 27752 30000 27872 0 FreeSans 480 0 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal3 s 29200 29792 30000 29912 0 FreeSans 480 0 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal3 s 29200 31832 30000 31952 0 FreeSans 480 0 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 27066 33200 27122 34000 0 FreeSans 224 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 23754 33200 23810 34000 0 FreeSans 224 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 20442 33200 20498 34000 0 FreeSans 224 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 17130 33200 17186 34000 0 FreeSans 224 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 13818 33200 13874 34000 0 FreeSans 224 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal3 s 29200 5312 30000 5432 0 FreeSans 480 0 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 10506 33200 10562 34000 0 FreeSans 224 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 7194 33200 7250 34000 0 FreeSans 224 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 3882 33200 3938 34000 0 FreeSans 224 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 570 33200 626 34000 0 FreeSans 224 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s 0 29520 800 29640 0 FreeSans 480 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal3 s 0 27480 800 27600 0 FreeSans 480 0 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal3 s 0 25440 800 25560 0 FreeSans 480 0 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal3 s 0 23400 800 23520 0 FreeSans 480 0 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s 0 21360 800 21480 0 FreeSans 480 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal3 s 0 19320 800 19440 0 FreeSans 480 0 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal3 s 29200 7352 30000 7472 0 FreeSans 480 0 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal3 s 0 17280 800 17400 0 FreeSans 480 0 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s 0 15240 800 15360 0 FreeSans 480 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal3 s 0 13200 800 13320 0 FreeSans 480 0 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s 0 9120 800 9240 0 FreeSans 480 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal3 s 0 7080 800 7200 0 FreeSans 480 0 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal3 s 0 5040 800 5160 0 FreeSans 480 0 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s 0 3000 800 3120 0 FreeSans 480 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 29200 9392 30000 9512 0 FreeSans 480 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal3 s 29200 11432 30000 11552 0 FreeSans 480 0 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal3 s 29200 13472 30000 13592 0 FreeSans 480 0 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal3 s 29200 15512 30000 15632 0 FreeSans 480 0 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal3 s 29200 17552 30000 17672 0 FreeSans 480 0 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 29200 19592 30000 19712 0 FreeSans 480 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal3 s 29200 21632 30000 21752 0 FreeSans 480 0 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 29200 2592 30000 2712 0 FreeSans 480 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal3 s 29200 22992 30000 23112 0 FreeSans 480 0 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 29200 25032 30000 25152 0 FreeSans 480 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 29200 27072 30000 27192 0 FreeSans 480 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 29200 29112 30000 29232 0 FreeSans 480 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal3 s 29200 31152 30000 31272 0 FreeSans 480 0 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 28170 33200 28226 34000 0 FreeSans 224 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 24858 33200 24914 34000 0 FreeSans 224 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 21546 33200 21602 34000 0 FreeSans 224 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 18234 33200 18290 34000 0 FreeSans 224 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 14922 33200 14978 34000 0 FreeSans 224 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal3 s 29200 4632 30000 4752 0 FreeSans 480 0 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 11610 33200 11666 34000 0 FreeSans 224 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 8298 33200 8354 34000 0 FreeSans 224 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 4986 33200 5042 34000 0 FreeSans 224 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 1674 33200 1730 34000 0 FreeSans 224 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal3 s 0 30200 800 30320 0 FreeSans 480 0 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal3 s 0 28160 800 28280 0 FreeSans 480 0 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal3 s 0 26120 800 26240 0 FreeSans 480 0 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal3 s 0 24080 800 24200 0 FreeSans 480 0 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal3 s 0 22040 800 22160 0 FreeSans 480 0 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal3 s 0 20000 800 20120 0 FreeSans 480 0 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 29200 6672 30000 6792 0 FreeSans 480 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s 0 17960 800 18080 0 FreeSans 480 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal3 s 0 15920 800 16040 0 FreeSans 480 0 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal3 s 0 13880 800 14000 0 FreeSans 480 0 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal3 s 0 11840 800 11960 0 FreeSans 480 0 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s 0 9800 800 9920 0 FreeSans 480 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal3 s 0 7760 800 7880 0 FreeSans 480 0 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal3 s 0 5720 800 5840 0 FreeSans 480 0 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal3 s 0 3680 800 3800 0 FreeSans 480 0 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal3 s 29200 8712 30000 8832 0 FreeSans 480 0 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal3 s 29200 10752 30000 10872 0 FreeSans 480 0 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal3 s 29200 12792 30000 12912 0 FreeSans 480 0 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal3 s 29200 14832 30000 14952 0 FreeSans 480 0 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 29200 16872 30000 16992 0 FreeSans 480 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal3 s 29200 18912 30000 19032 0 FreeSans 480 0 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 29200 20952 30000 21072 0 FreeSans 480 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal4 s 4417 2128 4737 31600 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 11363 2128 11683 31600 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 18309 2128 18629 31600 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 25255 2128 25575 31600 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 7890 2128 8210 31600 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
flabel metal4 s 14836 2128 15156 31600 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
flabel metal4 s 21782 2128 22102 31600 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
flabel metal4 s 28728 2128 29048 31600 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
rlabel metal1 14996 31008 14996 31008 0 vccd1
rlabel via1 15076 31552 15076 31552 0 vssd1
rlabel metal1 16008 27914 16008 27914 0 _000_
rlabel metal1 5980 25398 5980 25398 0 _001_
rlabel metal1 16376 29274 16376 29274 0 _002_
rlabel metal2 10626 28560 10626 28560 0 _003_
rlabel metal1 15456 28730 15456 28730 0 _004_
rlabel metal1 10856 24378 10856 24378 0 _005_
rlabel metal1 9614 29580 9614 29580 0 _006_
rlabel metal1 2548 31382 2548 31382 0 _007_
rlabel metal1 8648 23834 8648 23834 0 _008_
rlabel metal1 2323 30090 2323 30090 0 _009_
rlabel metal1 8004 25398 8004 25398 0 _010_
rlabel metal3 13340 27472 13340 27472 0 _011_
rlabel metal2 3450 28424 3450 28424 0 _012_
rlabel metal2 18722 30481 18722 30481 0 _013_
rlabel metal2 12742 30243 12742 30243 0 _014_
rlabel metal1 14781 30294 14781 30294 0 _015_
rlabel metal1 16560 27574 16560 27574 0 _016_
rlabel via2 11730 25925 11730 25925 0 _017_
rlabel via2 2622 29563 2622 29563 0 _018_
rlabel metal1 12047 28050 12047 28050 0 _019_
rlabel metal2 3266 26741 3266 26741 0 _020_
rlabel metal1 9839 28118 9839 28118 0 _021_
rlabel metal2 15318 29920 15318 29920 0 _022_
rlabel via2 19826 30821 19826 30821 0 _023_
rlabel metal1 12972 27098 12972 27098 0 _024_
rlabel metal1 5612 26486 5612 26486 0 _025_
rlabel metal1 6578 26486 6578 26486 0 _026_
rlabel metal1 8786 25466 8786 25466 0 _027_
rlabel metal1 4646 27642 4646 27642 0 _028_
rlabel metal2 2346 29699 2346 29699 0 _029_
rlabel metal1 5336 27098 5336 27098 0 _030_
rlabel metal1 9292 27030 9292 27030 0 _031_
rlabel metal2 15962 28322 15962 28322 0 _032_
rlabel metal1 16100 27846 16100 27846 0 _033_
rlabel metal1 17618 28730 17618 28730 0 _034_
rlabel metal1 17066 28458 17066 28458 0 _035_
rlabel metal2 10350 26027 10350 26027 0 _036_
rlabel metal1 19366 30124 19366 30124 0 _037_
rlabel metal1 17158 30260 17158 30260 0 _038_
rlabel metal2 16882 26588 16882 26588 0 _039_
rlabel metal2 16698 25874 16698 25874 0 _040_
rlabel metal1 13616 27506 13616 27506 0 _041_
rlabel metal2 13202 26044 13202 26044 0 _042_
rlabel metal1 12834 27506 12834 27506 0 _043_
rlabel metal1 15318 27846 15318 27846 0 _044_
rlabel via2 13202 27421 13202 27421 0 _045_
rlabel via2 15042 28067 15042 28067 0 _046_
rlabel metal1 7314 25738 7314 25738 0 _047_
rlabel metal2 12650 25432 12650 25432 0 _048_
rlabel metal1 12696 26894 12696 26894 0 _049_
rlabel metal1 13616 25874 13616 25874 0 _050_
rlabel metal1 15548 25670 15548 25670 0 _051_
rlabel metal1 15456 29614 15456 29614 0 _052_
rlabel metal2 16882 29886 16882 29886 0 _053_
rlabel metal2 15134 27404 15134 27404 0 _054_
rlabel metal3 13570 28492 13570 28492 0 _055_
rlabel metal1 2254 26384 2254 26384 0 _056_
rlabel via2 13202 26979 13202 26979 0 _057_
rlabel metal1 5750 26384 5750 26384 0 _058_
rlabel metal1 6072 25738 6072 25738 0 _059_
rlabel metal1 4876 29614 4876 29614 0 _060_
rlabel metal1 6394 26350 6394 26350 0 _061_
rlabel metal1 7406 24174 7406 24174 0 _062_
rlabel metal2 8418 24820 8418 24820 0 _063_
rlabel metal2 1978 29308 1978 29308 0 _064_
rlabel metal1 5796 24650 5796 24650 0 _065_
rlabel metal2 2162 27438 2162 27438 0 _066_
rlabel metal1 3956 26962 3956 26962 0 _067_
rlabel metal1 4140 26962 4140 26962 0 _068_
rlabel metal2 6578 31484 6578 31484 0 _069_
rlabel metal2 13846 26078 13846 26078 0 _070_
rlabel metal1 20286 30770 20286 30770 0 _071_
rlabel metal1 16238 30906 16238 30906 0 _072_
rlabel via2 13662 26435 13662 26435 0 _073_
rlabel metal1 15962 28730 15962 28730 0 _074_
rlabel metal2 2714 25500 2714 25500 0 _075_
rlabel metal1 20532 31382 20532 31382 0 _076_
rlabel metal2 13294 30702 13294 30702 0 _077_
rlabel metal1 12558 25296 12558 25296 0 _078_
rlabel metal2 10810 24378 10810 24378 0 _079_
rlabel metal1 17940 30226 17940 30226 0 _080_
rlabel metal2 20286 30192 20286 30192 0 _081_
rlabel metal1 17572 29138 17572 29138 0 _082_
rlabel metal1 12742 26282 12742 26282 0 _083_
rlabel metal2 10626 25177 10626 25177 0 _084_
rlabel metal1 6394 29138 6394 29138 0 _085_
rlabel metal1 2622 30192 2622 30192 0 _086_
rlabel metal1 9200 23698 9200 23698 0 _087_
rlabel metal2 2070 29087 2070 29087 0 _088_
rlabel metal1 5152 25330 5152 25330 0 _089_
rlabel metal1 7590 25228 7590 25228 0 _090_
rlabel metal1 14904 26826 14904 26826 0 _091_
rlabel metal2 11730 24735 11730 24735 0 _092_
rlabel metal1 11868 28730 11868 28730 0 clknet_0_io_in[0]
rlabel metal1 7682 29614 7682 29614 0 clknet_2_0__leaf_io_in[0]
rlabel metal2 2714 29682 2714 29682 0 clknet_2_1__leaf_io_in[0]
rlabel metal1 11224 27506 11224 27506 0 clknet_2_2__leaf_io_in[0]
rlabel metal1 12282 30838 12282 30838 0 clknet_2_3__leaf_io_in[0]
rlabel metal3 12719 27948 12719 27948 0 io_in[0]
rlabel via2 28382 4029 28382 4029 0 io_in[1]
rlabel metal1 18538 30090 18538 30090 0 io_out[18]
rlabel metal1 12512 29274 12512 29274 0 io_out[19]
rlabel metal2 11822 33252 11822 33252 0 io_out[20]
rlabel metal1 7728 24650 7728 24650 0 io_out[21]
rlabel metal1 4922 26554 4922 26554 0 io_out[22]
rlabel metal1 2116 26826 2116 26826 0 io_out[23]
rlabel metal2 2898 28679 2898 28679 0 io_out[24]
rlabel metal3 1188 28220 1188 28220 0 io_out[25]
rlabel via2 7038 30277 7038 30277 0 mod._autorun
rlabel metal1 15686 27370 15686 27370 0 mod._d_io_out\[0\]
rlabel metal1 12926 26928 12926 26928 0 mod._d_io_out\[1\]
rlabel metal1 6026 25874 6026 25874 0 mod._d_io_out\[2\]
rlabel metal1 5842 25942 5842 25942 0 mod._d_io_out\[3\]
rlabel metal1 4646 29546 4646 29546 0 mod._d_io_out\[4\]
rlabel metal1 4922 29784 4922 29784 0 mod._d_io_out\[5\]
rlabel metal1 1886 29036 1886 29036 0 mod._d_io_out\[6\]
rlabel metal1 7728 26350 7728 26350 0 mod._d_io_out\[7\]
rlabel metal2 19734 30940 19734 30940 0 mod._q_cnt\[0\]
rlabel metal2 15870 28254 15870 28254 0 mod._q_cnt\[10\]
rlabel metal1 13386 30600 13386 30600 0 mod._q_cnt\[11\]
rlabel metal1 14306 30022 14306 30022 0 mod._q_cnt\[12\]
rlabel metal2 9890 25500 9890 25500 0 mod._q_cnt\[13\]
rlabel metal2 6026 29223 6026 29223 0 mod._q_cnt\[14\]
rlabel metal2 13478 27353 13478 27353 0 mod._q_cnt\[15\]
rlabel metal1 15916 27982 15916 27982 0 mod._q_cnt\[16\]
rlabel metal2 13018 25993 13018 25993 0 mod._q_cnt\[17\]
rlabel metal3 14858 28900 14858 28900 0 mod._q_cnt\[18\]
rlabel metal2 14582 30005 14582 30005 0 mod._q_cnt\[19\]
rlabel metal2 11362 31280 11362 31280 0 mod._q_cnt\[1\]
rlabel metal2 19642 30702 19642 30702 0 mod._q_cnt\[2\]
rlabel metal2 16698 30345 16698 30345 0 mod._q_cnt\[3\]
rlabel metal2 8418 30736 8418 30736 0 mod._q_cnt\[4\]
rlabel metal1 8556 26350 8556 26350 0 mod._q_cnt\[5\]
rlabel metal1 2346 30260 2346 30260 0 mod._q_cnt\[6\]
rlabel metal2 8418 27200 8418 27200 0 mod._q_cnt\[7\]
rlabel metal2 14398 27778 14398 27778 0 mod._q_cnt\[8\]
rlabel metal2 8418 26826 8418 26826 0 mod._q_cnt\[9\]
rlabel metal1 19036 30566 19036 30566 0 mod._q_index\[0\]
rlabel metal1 11776 29750 11776 29750 0 mod._q_index\[1\]
rlabel metal1 17388 25874 17388 25874 0 net1
rlabel metal3 1142 3060 1142 3060 0 net10
rlabel metal3 28850 2652 28850 2652 0 net11
rlabel metal2 28382 4845 28382 4845 0 net12
rlabel via2 28382 6749 28382 6749 0 net13
rlabel via2 28382 9061 28382 9061 0 net14
rlabel via2 28382 11101 28382 11101 0 net15
rlabel metal2 28382 13073 28382 13073 0 net16
rlabel via2 28382 14875 28382 14875 0 net17
rlabel via2 28382 16949 28382 16949 0 net18
rlabel metal2 28382 19057 28382 19057 0 net19
rlabel metal1 18400 30226 18400 30226 0 net2
rlabel metal2 28382 21165 28382 21165 0 net20
rlabel via2 28382 23069 28382 23069 0 net21
rlabel via2 28382 25381 28382 25381 0 net22
rlabel via2 28382 27421 28382 27421 0 net23
rlabel metal2 28382 29393 28382 29393 0 net24
rlabel metal2 28382 31059 28382 31059 0 net25
rlabel metal2 28198 32276 28198 32276 0 net26
rlabel metal1 24932 31314 24932 31314 0 net27
rlabel metal1 21804 31314 21804 31314 0 net28
rlabel metal3 1142 26180 1142 26180 0 net29
rlabel metal1 11776 29138 11776 29138 0 net3
rlabel metal3 1142 24140 1142 24140 0 net30
rlabel metal3 1142 22100 1142 22100 0 net31
rlabel metal3 1142 20060 1142 20060 0 net32
rlabel metal3 1142 18020 1142 18020 0 net33
rlabel metal3 1142 15980 1142 15980 0 net34
rlabel metal3 1142 13940 1142 13940 0 net35
rlabel metal3 1142 11900 1142 11900 0 net36
rlabel metal3 1142 9860 1142 9860 0 net37
rlabel metal3 1142 7820 1142 7820 0 net38
rlabel metal3 1142 5780 1142 5780 0 net39
rlabel metal1 11178 29580 11178 29580 0 net4
rlabel metal3 1142 3740 1142 3740 0 net40
rlabel via2 28382 3621 28382 3621 0 net41
rlabel via2 28382 5661 28382 5661 0 net42
rlabel metal2 28382 7633 28382 7633 0 net43
rlabel via2 28382 9435 28382 9435 0 net44
rlabel via2 28382 11509 28382 11509 0 net45
rlabel metal2 28382 13617 28382 13617 0 net46
rlabel metal2 28382 15725 28382 15725 0 net47
rlabel via2 28382 17629 28382 17629 0 net48
rlabel via2 28382 19941 28382 19941 0 net49
rlabel metal1 7498 24752 7498 24752 0 net5
rlabel via2 28382 21981 28382 21981 0 net50
rlabel metal2 28382 23953 28382 23953 0 net51
rlabel via2 28382 25755 28382 25755 0 net52
rlabel via2 28382 27829 28382 27829 0 net53
rlabel metal2 28382 29937 28382 29937 0 net54
rlabel metal3 28528 31892 28528 31892 0 net55
rlabel metal1 27140 31314 27140 31314 0 net56
rlabel metal1 23828 31314 23828 31314 0 net57
rlabel metal2 20470 32489 20470 32489 0 net58
rlabel metal2 17158 32489 17158 32489 0 net59
rlabel metal1 4508 26350 4508 26350 0 net6
rlabel metal2 16146 31586 16146 31586 0 net60
rlabel metal2 10718 33252 10718 33252 0 net61
rlabel metal2 7038 33252 7038 33252 0 net62
rlabel metal1 3956 25874 3956 25874 0 net63
rlabel metal2 276 33252 276 33252 0 net64
rlabel metal3 1119 29580 1119 29580 0 net65
rlabel metal2 2806 26469 2806 26469 0 net66
rlabel metal3 1510 25500 1510 25500 0 net67
rlabel metal3 1142 23460 1142 23460 0 net68
rlabel metal3 1142 21420 1142 21420 0 net69
rlabel metal1 2622 26894 2622 26894 0 net7
rlabel metal3 1142 19380 1142 19380 0 net70
rlabel metal3 1142 17340 1142 17340 0 net71
rlabel metal3 1142 15300 1142 15300 0 net72
rlabel metal3 1142 13260 1142 13260 0 net73
rlabel metal3 1142 11220 1142 11220 0 net74
rlabel metal3 1142 9180 1142 9180 0 net75
rlabel metal3 1142 7140 1142 7140 0 net76
rlabel metal3 1142 5100 1142 5100 0 net77
rlabel metal2 7222 26792 7222 26792 0 net78
rlabel metal1 3261 28458 3261 28458 0 net79
rlabel metal1 1886 26996 1886 26996 0 net8
rlabel metal1 1886 25908 1886 25908 0 net9
<< properties >>
string FIXED_BBOX 0 0 30000 34000
<< end >>
