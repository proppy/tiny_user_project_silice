// This is the unpowered netlist.
module tiny_user_project (io_in,
    io_oeb,
    io_out);
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire net42;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net43;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net44;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net11;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net12;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net13;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net14;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire \mod._autorun ;
 wire \mod._d_io_out[0] ;
 wire \mod._d_io_out[1] ;
 wire \mod._d_io_out[2] ;
 wire \mod._d_io_out[3] ;
 wire \mod._d_io_out[4] ;
 wire \mod._d_io_out[5] ;
 wire \mod._d_io_out[6] ;
 wire \mod._d_io_out[7] ;
 wire \mod._q_cnt[0] ;
 wire \mod._q_cnt[10] ;
 wire \mod._q_cnt[11] ;
 wire \mod._q_cnt[12] ;
 wire \mod._q_cnt[13] ;
 wire \mod._q_cnt[14] ;
 wire \mod._q_cnt[15] ;
 wire \mod._q_cnt[16] ;
 wire \mod._q_cnt[17] ;
 wire \mod._q_cnt[18] ;
 wire \mod._q_cnt[19] ;
 wire \mod._q_cnt[1] ;
 wire \mod._q_cnt[2] ;
 wire \mod._q_cnt[3] ;
 wire \mod._q_cnt[4] ;
 wire \mod._q_cnt[5] ;
 wire \mod._q_cnt[6] ;
 wire \mod._q_cnt[7] ;
 wire \mod._q_cnt[8] ;
 wire \mod._q_cnt[9] ;
 wire \mod._q_index[0] ;
 wire \mod._q_index[1] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net78;
 wire net79;
 wire [0:0] clknet_0_io_in;
 wire [0:0] clknet_2_0__leaf_io_in;
 wire [0:0] clknet_2_1__leaf_io_in;
 wire [0:0] clknet_2_2__leaf_io_in;
 wire [0:0] clknet_2_3__leaf_io_in;

 sky130_fd_sc_hd__buf_2 _093_ (.A(net1),
    .X(_069_));
 sky130_fd_sc_hd__inv_2 _094_ (.A(_069_),
    .Y(_000_));
 sky130_fd_sc_hd__or2_1 _095_ (.A(\mod._autorun ),
    .B(_069_),
    .X(_070_));
 sky130_fd_sc_hd__clkbuf_1 _096_ (.A(_070_),
    .X(_001_));
 sky130_fd_sc_hd__clkbuf_2 _097_ (.A(_069_),
    .X(_071_));
 sky130_fd_sc_hd__a21o_1 _098_ (.A1(\mod._q_index[1] ),
    .A2(\mod._autorun ),
    .B1(_071_),
    .X(_002_));
 sky130_fd_sc_hd__inv_2 _099_ (.A(\mod._q_index[1] ),
    .Y(_072_));
 sky130_fd_sc_hd__a21oi_1 _100_ (.A1(_072_),
    .A2(\mod._q_index[0] ),
    .B1(\mod._q_cnt[0] ),
    .Y(_073_));
 sky130_fd_sc_hd__and3_1 _101_ (.A(\mod._q_cnt[0] ),
    .B(_072_),
    .C(\mod._q_index[0] ),
    .X(_074_));
 sky130_fd_sc_hd__nor3_1 _102_ (.A(_071_),
    .B(_073_),
    .C(_074_),
    .Y(_003_));
 sky130_fd_sc_hd__clkbuf_2 _103_ (.A(_069_),
    .X(_075_));
 sky130_fd_sc_hd__and4b_1 _104_ (.A_N(\mod._q_index[1] ),
    .B(\mod._q_index[0] ),
    .C(\mod._q_cnt[1] ),
    .D(\mod._q_cnt[0] ),
    .X(_076_));
 sky130_fd_sc_hd__nor2_1 _105_ (.A(_075_),
    .B(_076_),
    .Y(_077_));
 sky130_fd_sc_hd__o21a_1 _106_ (.A1(\mod._q_cnt[1] ),
    .A2(_074_),
    .B1(_077_),
    .X(_004_));
 sky130_fd_sc_hd__and2_1 _107_ (.A(\mod._q_cnt[2] ),
    .B(_076_),
    .X(_078_));
 sky130_fd_sc_hd__o21ai_1 _108_ (.A1(\mod._q_cnt[2] ),
    .A2(_076_),
    .B1(_000_),
    .Y(_079_));
 sky130_fd_sc_hd__nor2_1 _109_ (.A(_078_),
    .B(_079_),
    .Y(_005_));
 sky130_fd_sc_hd__and3_1 _110_ (.A(\mod._q_cnt[3] ),
    .B(\mod._q_cnt[2] ),
    .C(_076_),
    .X(_080_));
 sky130_fd_sc_hd__nor2_1 _111_ (.A(_075_),
    .B(_080_),
    .Y(_081_));
 sky130_fd_sc_hd__o21a_1 _112_ (.A1(\mod._q_cnt[3] ),
    .A2(_078_),
    .B1(_081_),
    .X(_006_));
 sky130_fd_sc_hd__and2_1 _113_ (.A(\mod._q_cnt[4] ),
    .B(_080_),
    .X(_082_));
 sky130_fd_sc_hd__nor2_1 _114_ (.A(_075_),
    .B(_082_),
    .Y(_083_));
 sky130_fd_sc_hd__o21a_1 _115_ (.A1(\mod._q_cnt[4] ),
    .A2(_080_),
    .B1(_083_),
    .X(_007_));
 sky130_fd_sc_hd__and2_1 _116_ (.A(\mod._q_cnt[5] ),
    .B(\mod._q_cnt[4] ),
    .X(_084_));
 sky130_fd_sc_hd__and4_1 _117_ (.A(\mod._q_cnt[3] ),
    .B(\mod._q_cnt[2] ),
    .C(_076_),
    .D(_084_),
    .X(_085_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _118_ (.A(_085_),
    .X(_086_));
 sky130_fd_sc_hd__o21ai_1 _119_ (.A1(\mod._q_cnt[5] ),
    .A2(_082_),
    .B1(_000_),
    .Y(_087_));
 sky130_fd_sc_hd__nor2_1 _120_ (.A(_086_),
    .B(_087_),
    .Y(_008_));
 sky130_fd_sc_hd__a21oi_1 _121_ (.A1(\mod._q_cnt[6] ),
    .A2(_086_),
    .B1(_071_),
    .Y(_088_));
 sky130_fd_sc_hd__o21a_1 _122_ (.A1(\mod._q_cnt[6] ),
    .A2(_086_),
    .B1(_088_),
    .X(_009_));
 sky130_fd_sc_hd__a21oi_1 _123_ (.A1(\mod._q_cnt[6] ),
    .A2(_086_),
    .B1(\mod._q_cnt[7] ),
    .Y(_089_));
 sky130_fd_sc_hd__and3_1 _124_ (.A(\mod._q_cnt[7] ),
    .B(\mod._q_cnt[6] ),
    .C(_086_),
    .X(_090_));
 sky130_fd_sc_hd__nor3_1 _125_ (.A(_071_),
    .B(_089_),
    .C(_090_),
    .Y(_010_));
 sky130_fd_sc_hd__a21oi_1 _126_ (.A1(\mod._q_cnt[8] ),
    .A2(_090_),
    .B1(_071_),
    .Y(_091_));
 sky130_fd_sc_hd__o21a_1 _127_ (.A1(\mod._q_cnt[8] ),
    .A2(_090_),
    .B1(_091_),
    .X(_011_));
 sky130_fd_sc_hd__a21oi_1 _128_ (.A1(\mod._q_cnt[8] ),
    .A2(_090_),
    .B1(\mod._q_cnt[9] ),
    .Y(_092_));
 sky130_fd_sc_hd__and2_1 _129_ (.A(\mod._q_cnt[9] ),
    .B(\mod._q_cnt[8] ),
    .X(_031_));
 sky130_fd_sc_hd__and4_1 _130_ (.A(\mod._q_cnt[7] ),
    .B(\mod._q_cnt[6] ),
    .C(_086_),
    .D(_031_),
    .X(_032_));
 sky130_fd_sc_hd__nor3_1 _131_ (.A(_071_),
    .B(_092_),
    .C(_032_),
    .Y(_012_));
 sky130_fd_sc_hd__and2_1 _132_ (.A(\mod._q_cnt[10] ),
    .B(_032_),
    .X(_033_));
 sky130_fd_sc_hd__o21ai_1 _133_ (.A1(\mod._q_cnt[10] ),
    .A2(_032_),
    .B1(_000_),
    .Y(_034_));
 sky130_fd_sc_hd__nor2_1 _134_ (.A(_033_),
    .B(_034_),
    .Y(_013_));
 sky130_fd_sc_hd__and3_1 _135_ (.A(\mod._q_cnt[11] ),
    .B(\mod._q_cnt[10] ),
    .C(_032_),
    .X(_035_));
 sky130_fd_sc_hd__nor2_1 _136_ (.A(_075_),
    .B(_035_),
    .Y(_036_));
 sky130_fd_sc_hd__o21a_1 _137_ (.A1(\mod._q_cnt[11] ),
    .A2(_033_),
    .B1(_036_),
    .X(_014_));
 sky130_fd_sc_hd__and4_1 _138_ (.A(\mod._q_cnt[12] ),
    .B(\mod._q_cnt[11] ),
    .C(\mod._q_cnt[10] ),
    .D(_032_),
    .X(_037_));
 sky130_fd_sc_hd__nor2_1 _139_ (.A(_075_),
    .B(_037_),
    .Y(_038_));
 sky130_fd_sc_hd__o21a_1 _140_ (.A1(\mod._q_cnt[12] ),
    .A2(_035_),
    .B1(_038_),
    .X(_015_));
 sky130_fd_sc_hd__and2_1 _141_ (.A(\mod._q_cnt[13] ),
    .B(_037_),
    .X(_039_));
 sky130_fd_sc_hd__o21ai_1 _142_ (.A1(\mod._q_cnt[13] ),
    .A2(_037_),
    .B1(_000_),
    .Y(_040_));
 sky130_fd_sc_hd__nor2_1 _143_ (.A(_039_),
    .B(_040_),
    .Y(_016_));
 sky130_fd_sc_hd__and3_1 _144_ (.A(\mod._q_cnt[14] ),
    .B(\mod._q_cnt[13] ),
    .C(_037_),
    .X(_041_));
 sky130_fd_sc_hd__nor2_1 _145_ (.A(_075_),
    .B(_041_),
    .Y(_042_));
 sky130_fd_sc_hd__o21a_1 _146_ (.A1(\mod._q_cnt[14] ),
    .A2(_039_),
    .B1(_042_),
    .X(_017_));
 sky130_fd_sc_hd__and4_1 _147_ (.A(\mod._q_cnt[15] ),
    .B(\mod._q_cnt[14] ),
    .C(\mod._q_cnt[13] ),
    .D(_037_),
    .X(_043_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _148_ (.A(_043_),
    .X(_044_));
 sky130_fd_sc_hd__nor2_1 _149_ (.A(_075_),
    .B(_044_),
    .Y(_045_));
 sky130_fd_sc_hd__o21a_1 _150_ (.A1(\mod._q_cnt[15] ),
    .A2(_041_),
    .B1(_045_),
    .X(_018_));
 sky130_fd_sc_hd__a21oi_1 _151_ (.A1(\mod._q_cnt[16] ),
    .A2(_044_),
    .B1(_071_),
    .Y(_046_));
 sky130_fd_sc_hd__o21a_1 _152_ (.A1(\mod._q_cnt[16] ),
    .A2(_044_),
    .B1(_046_),
    .X(_019_));
 sky130_fd_sc_hd__a21oi_1 _153_ (.A1(\mod._q_cnt[16] ),
    .A2(_044_),
    .B1(\mod._q_cnt[17] ),
    .Y(_047_));
 sky130_fd_sc_hd__and3_1 _154_ (.A(\mod._q_cnt[17] ),
    .B(\mod._q_cnt[16] ),
    .C(_044_),
    .X(_048_));
 sky130_fd_sc_hd__nor3_1 _155_ (.A(_071_),
    .B(_047_),
    .C(_048_),
    .Y(_020_));
 sky130_fd_sc_hd__and4_1 _156_ (.A(\mod._q_cnt[18] ),
    .B(\mod._q_cnt[17] ),
    .C(\mod._q_cnt[16] ),
    .D(_044_),
    .X(_049_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _157_ (.A(_049_),
    .X(_050_));
 sky130_fd_sc_hd__nor2_1 _158_ (.A(_069_),
    .B(_050_),
    .Y(_051_));
 sky130_fd_sc_hd__o21a_1 _159_ (.A1(\mod._q_cnt[18] ),
    .A2(_048_),
    .B1(_051_),
    .X(_021_));
 sky130_fd_sc_hd__a21oi_1 _160_ (.A1(\mod._q_cnt[19] ),
    .A2(_050_),
    .B1(_075_),
    .Y(_052_));
 sky130_fd_sc_hd__o21a_1 _161_ (.A1(\mod._q_cnt[19] ),
    .A2(_050_),
    .B1(_052_),
    .X(_022_));
 sky130_fd_sc_hd__a21oi_1 _162_ (.A1(\mod._q_cnt[19] ),
    .A2(_050_),
    .B1(\mod._d_io_out[0] ),
    .Y(_053_));
 sky130_fd_sc_hd__and3_1 _163_ (.A(\mod._d_io_out[0] ),
    .B(\mod._q_cnt[19] ),
    .C(_050_),
    .X(_054_));
 sky130_fd_sc_hd__nor3_1 _164_ (.A(_071_),
    .B(_053_),
    .C(_054_),
    .Y(_023_));
 sky130_fd_sc_hd__and4_1 _165_ (.A(\mod._d_io_out[1] ),
    .B(\mod._d_io_out[0] ),
    .C(\mod._q_cnt[19] ),
    .D(_050_),
    .X(_055_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _166_ (.A(_055_),
    .X(_056_));
 sky130_fd_sc_hd__nor2_1 _167_ (.A(_069_),
    .B(_056_),
    .Y(_057_));
 sky130_fd_sc_hd__o21a_1 _168_ (.A1(\mod._d_io_out[1] ),
    .A2(_054_),
    .B1(_057_),
    .X(_024_));
 sky130_fd_sc_hd__a21oi_1 _169_ (.A1(\mod._d_io_out[2] ),
    .A2(_056_),
    .B1(_075_),
    .Y(_058_));
 sky130_fd_sc_hd__o21a_1 _170_ (.A1(\mod._d_io_out[2] ),
    .A2(_056_),
    .B1(_058_),
    .X(_025_));
 sky130_fd_sc_hd__a21oi_1 _171_ (.A1(\mod._d_io_out[2] ),
    .A2(_056_),
    .B1(\mod._d_io_out[3] ),
    .Y(_059_));
 sky130_fd_sc_hd__and2_1 _172_ (.A(\mod._d_io_out[3] ),
    .B(\mod._d_io_out[2] ),
    .X(_060_));
 sky130_fd_sc_hd__and2_1 _173_ (.A(_056_),
    .B(_060_),
    .X(_061_));
 sky130_fd_sc_hd__nor3_1 _174_ (.A(_071_),
    .B(_059_),
    .C(_061_),
    .Y(_026_));
 sky130_fd_sc_hd__and3_1 _175_ (.A(\mod._d_io_out[4] ),
    .B(_056_),
    .C(_060_),
    .X(_062_));
 sky130_fd_sc_hd__nor2_1 _176_ (.A(_069_),
    .B(_062_),
    .Y(_063_));
 sky130_fd_sc_hd__o21a_1 _177_ (.A1(\mod._d_io_out[4] ),
    .A2(_061_),
    .B1(_063_),
    .X(_027_));
 sky130_fd_sc_hd__and4_1 _178_ (.A(\mod._d_io_out[5] ),
    .B(\mod._d_io_out[4] ),
    .C(_056_),
    .D(_060_),
    .X(_064_));
 sky130_fd_sc_hd__nor2_1 _179_ (.A(_069_),
    .B(_064_),
    .Y(_065_));
 sky130_fd_sc_hd__o21a_1 _180_ (.A1(\mod._d_io_out[5] ),
    .A2(_062_),
    .B1(_065_),
    .X(_028_));
 sky130_fd_sc_hd__a21oi_1 _181_ (.A1(\mod._d_io_out[6] ),
    .A2(_064_),
    .B1(_075_),
    .Y(_066_));
 sky130_fd_sc_hd__o21a_1 _182_ (.A1(\mod._d_io_out[6] ),
    .A2(_064_),
    .B1(_066_),
    .X(_029_));
 sky130_fd_sc_hd__a21oi_1 _183_ (.A1(\mod._d_io_out[6] ),
    .A2(_064_),
    .B1(\mod._d_io_out[7] ),
    .Y(_067_));
 sky130_fd_sc_hd__a31o_1 _184_ (.A1(\mod._d_io_out[7] ),
    .A2(\mod._d_io_out[6] ),
    .A3(_064_),
    .B1(_069_),
    .X(_068_));
 sky130_fd_sc_hd__nor2_1 _185_ (.A(_067_),
    .B(_068_),
    .Y(_030_));
 sky130_fd_sc_hd__dfxtp_1 _186_ (.CLK(clknet_2_1__leaf_io_in[0]),
    .D(_000_),
    .Q(\mod._autorun ));
 sky130_fd_sc_hd__dfxtp_1 _187_ (.CLK(clknet_2_1__leaf_io_in[0]),
    .D(_001_),
    .Q(\mod._q_index[0] ));
 sky130_fd_sc_hd__dfxtp_1 _188_ (.CLK(clknet_2_3__leaf_io_in[0]),
    .D(_002_),
    .Q(\mod._q_index[1] ));
 sky130_fd_sc_hd__dfxtp_1 _189_ (.CLK(clknet_2_3__leaf_io_in[0]),
    .D(\mod._d_io_out[0] ),
    .Q(net2));
 sky130_fd_sc_hd__dfxtp_1 _190_ (.CLK(clknet_2_3__leaf_io_in[0]),
    .D(\mod._d_io_out[1] ),
    .Q(net3));
 sky130_fd_sc_hd__dfxtp_1 _191_ (.CLK(clknet_2_2__leaf_io_in[0]),
    .D(\mod._d_io_out[2] ),
    .Q(net4));
 sky130_fd_sc_hd__dfxtp_1 _192_ (.CLK(clknet_2_1__leaf_io_in[0]),
    .D(net79),
    .Q(net5));
 sky130_fd_sc_hd__dfxtp_1 _193_ (.CLK(clknet_2_1__leaf_io_in[0]),
    .D(\mod._d_io_out[4] ),
    .Q(net6));
 sky130_fd_sc_hd__dfxtp_1 _194_ (.CLK(clknet_2_0__leaf_io_in[0]),
    .D(\mod._d_io_out[5] ),
    .Q(net7));
 sky130_fd_sc_hd__dfxtp_1 _195_ (.CLK(clknet_2_1__leaf_io_in[0]),
    .D(\mod._d_io_out[6] ),
    .Q(net8));
 sky130_fd_sc_hd__dfxtp_1 _196_ (.CLK(clknet_2_1__leaf_io_in[0]),
    .D(net78),
    .Q(net9));
 sky130_fd_sc_hd__dfxtp_1 _197_ (.CLK(clknet_2_2__leaf_io_in[0]),
    .D(_003_),
    .Q(\mod._q_cnt[0] ));
 sky130_fd_sc_hd__dfxtp_1 _198_ (.CLK(clknet_2_1__leaf_io_in[0]),
    .D(_004_),
    .Q(\mod._q_cnt[1] ));
 sky130_fd_sc_hd__dfxtp_1 _199_ (.CLK(clknet_2_2__leaf_io_in[0]),
    .D(_005_),
    .Q(\mod._q_cnt[2] ));
 sky130_fd_sc_hd__dfxtp_1 _200_ (.CLK(clknet_2_0__leaf_io_in[0]),
    .D(_006_),
    .Q(\mod._q_cnt[3] ));
 sky130_fd_sc_hd__dfxtp_1 _201_ (.CLK(clknet_2_1__leaf_io_in[0]),
    .D(_007_),
    .Q(\mod._q_cnt[4] ));
 sky130_fd_sc_hd__dfxtp_1 _202_ (.CLK(clknet_2_0__leaf_io_in[0]),
    .D(_008_),
    .Q(\mod._q_cnt[5] ));
 sky130_fd_sc_hd__dfxtp_1 _203_ (.CLK(clknet_2_1__leaf_io_in[0]),
    .D(_009_),
    .Q(\mod._q_cnt[6] ));
 sky130_fd_sc_hd__dfxtp_1 _204_ (.CLK(clknet_2_0__leaf_io_in[0]),
    .D(_010_),
    .Q(\mod._q_cnt[7] ));
 sky130_fd_sc_hd__dfxtp_1 _205_ (.CLK(clknet_2_2__leaf_io_in[0]),
    .D(_011_),
    .Q(\mod._q_cnt[8] ));
 sky130_fd_sc_hd__dfxtp_1 _206_ (.CLK(clknet_2_0__leaf_io_in[0]),
    .D(_012_),
    .Q(\mod._q_cnt[9] ));
 sky130_fd_sc_hd__dfxtp_1 _207_ (.CLK(clknet_2_2__leaf_io_in[0]),
    .D(_013_),
    .Q(\mod._q_cnt[10] ));
 sky130_fd_sc_hd__dfxtp_1 _208_ (.CLK(clknet_2_3__leaf_io_in[0]),
    .D(_014_),
    .Q(\mod._q_cnt[11] ));
 sky130_fd_sc_hd__dfxtp_1 _209_ (.CLK(clknet_2_3__leaf_io_in[0]),
    .D(_015_),
    .Q(\mod._q_cnt[12] ));
 sky130_fd_sc_hd__dfxtp_1 _210_ (.CLK(clknet_2_3__leaf_io_in[0]),
    .D(_016_),
    .Q(\mod._q_cnt[13] ));
 sky130_fd_sc_hd__dfxtp_1 _211_ (.CLK(clknet_2_1__leaf_io_in[0]),
    .D(_017_),
    .Q(\mod._q_cnt[14] ));
 sky130_fd_sc_hd__dfxtp_1 _212_ (.CLK(clknet_2_1__leaf_io_in[0]),
    .D(_018_),
    .Q(\mod._q_cnt[15] ));
 sky130_fd_sc_hd__dfxtp_1 _213_ (.CLK(clknet_2_2__leaf_io_in[0]),
    .D(_019_),
    .Q(\mod._q_cnt[16] ));
 sky130_fd_sc_hd__dfxtp_1 _214_ (.CLK(clknet_2_0__leaf_io_in[0]),
    .D(_020_),
    .Q(\mod._q_cnt[17] ));
 sky130_fd_sc_hd__dfxtp_1 _215_ (.CLK(clknet_2_0__leaf_io_in[0]),
    .D(_021_),
    .Q(\mod._q_cnt[18] ));
 sky130_fd_sc_hd__dfxtp_1 _216_ (.CLK(clknet_2_3__leaf_io_in[0]),
    .D(_022_),
    .Q(\mod._q_cnt[19] ));
 sky130_fd_sc_hd__dfxtp_1 _217_ (.CLK(clknet_2_2__leaf_io_in[0]),
    .D(_023_),
    .Q(\mod._d_io_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 _218_ (.CLK(clknet_2_1__leaf_io_in[0]),
    .D(_024_),
    .Q(\mod._d_io_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 _219_ (.CLK(clknet_2_1__leaf_io_in[0]),
    .D(_025_),
    .Q(\mod._d_io_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 _220_ (.CLK(clknet_2_0__leaf_io_in[0]),
    .D(_026_),
    .Q(\mod._d_io_out[3] ));
 sky130_fd_sc_hd__dfxtp_1 _221_ (.CLK(clknet_2_0__leaf_io_in[0]),
    .D(_027_),
    .Q(\mod._d_io_out[4] ));
 sky130_fd_sc_hd__dfxtp_1 _222_ (.CLK(clknet_2_1__leaf_io_in[0]),
    .D(_028_),
    .Q(\mod._d_io_out[5] ));
 sky130_fd_sc_hd__dfxtp_1 _223_ (.CLK(clknet_2_3__leaf_io_in[0]),
    .D(_029_),
    .Q(\mod._d_io_out[6] ));
 sky130_fd_sc_hd__dfxtp_1 _224_ (.CLK(clknet_2_0__leaf_io_in[0]),
    .D(_030_),
    .Q(\mod._d_io_out[7] ));
 sky130_fd_sc_hd__conb_1 tiny_user_project_11 (.LO(net11));
 sky130_fd_sc_hd__conb_1 tiny_user_project_12 (.LO(net12));
 sky130_fd_sc_hd__conb_1 tiny_user_project_13 (.LO(net13));
 sky130_fd_sc_hd__conb_1 tiny_user_project_14 (.LO(net14));
 sky130_fd_sc_hd__conb_1 tiny_user_project_15 (.LO(net15));
 sky130_fd_sc_hd__conb_1 tiny_user_project_16 (.LO(net16));
 sky130_fd_sc_hd__conb_1 tiny_user_project_17 (.LO(net17));
 sky130_fd_sc_hd__conb_1 tiny_user_project_18 (.LO(net18));
 sky130_fd_sc_hd__conb_1 tiny_user_project_19 (.LO(net19));
 sky130_fd_sc_hd__conb_1 tiny_user_project_20 (.LO(net20));
 sky130_fd_sc_hd__conb_1 tiny_user_project_21 (.LO(net21));
 sky130_fd_sc_hd__conb_1 tiny_user_project_22 (.LO(net22));
 sky130_fd_sc_hd__conb_1 tiny_user_project_23 (.LO(net23));
 sky130_fd_sc_hd__conb_1 tiny_user_project_24 (.LO(net24));
 sky130_fd_sc_hd__conb_1 tiny_user_project_25 (.LO(net25));
 sky130_fd_sc_hd__conb_1 tiny_user_project_26 (.LO(net26));
 sky130_fd_sc_hd__conb_1 tiny_user_project_27 (.LO(net27));
 sky130_fd_sc_hd__conb_1 tiny_user_project_28 (.LO(net28));
 sky130_fd_sc_hd__conb_1 tiny_user_project_29 (.LO(net29));
 sky130_fd_sc_hd__conb_1 tiny_user_project_30 (.LO(net30));
 sky130_fd_sc_hd__conb_1 tiny_user_project_31 (.LO(net31));
 sky130_fd_sc_hd__conb_1 tiny_user_project_32 (.LO(net32));
 sky130_fd_sc_hd__conb_1 tiny_user_project_33 (.LO(net33));
 sky130_fd_sc_hd__conb_1 tiny_user_project_34 (.LO(net34));
 sky130_fd_sc_hd__conb_1 tiny_user_project_35 (.LO(net35));
 sky130_fd_sc_hd__conb_1 tiny_user_project_36 (.LO(net36));
 sky130_fd_sc_hd__conb_1 tiny_user_project_37 (.LO(net37));
 sky130_fd_sc_hd__conb_1 tiny_user_project_38 (.LO(net38));
 sky130_fd_sc_hd__conb_1 tiny_user_project_39 (.LO(net39));
 sky130_fd_sc_hd__conb_1 tiny_user_project_40 (.LO(net40));
 sky130_fd_sc_hd__conb_1 tiny_user_project_41 (.LO(net41));
 sky130_fd_sc_hd__conb_1 tiny_user_project_42 (.LO(net42));
 sky130_fd_sc_hd__conb_1 tiny_user_project_43 (.LO(net43));
 sky130_fd_sc_hd__conb_1 tiny_user_project_44 (.LO(net44));
 sky130_fd_sc_hd__conb_1 tiny_user_project_45 (.LO(net45));
 sky130_fd_sc_hd__conb_1 tiny_user_project_46 (.LO(net46));
 sky130_fd_sc_hd__conb_1 tiny_user_project_47 (.LO(net47));
 sky130_fd_sc_hd__conb_1 tiny_user_project_48 (.LO(net48));
 sky130_fd_sc_hd__conb_1 tiny_user_project_49 (.LO(net49));
 sky130_fd_sc_hd__conb_1 tiny_user_project_50 (.LO(net50));
 sky130_fd_sc_hd__conb_1 tiny_user_project_51 (.LO(net51));
 sky130_fd_sc_hd__conb_1 tiny_user_project_52 (.LO(net52));
 sky130_fd_sc_hd__conb_1 tiny_user_project_53 (.LO(net53));
 sky130_fd_sc_hd__conb_1 tiny_user_project_54 (.LO(net54));
 sky130_fd_sc_hd__conb_1 tiny_user_project_55 (.LO(net55));
 sky130_fd_sc_hd__conb_1 tiny_user_project_56 (.LO(net56));
 sky130_fd_sc_hd__conb_1 tiny_user_project_57 (.LO(net57));
 sky130_fd_sc_hd__conb_1 tiny_user_project_58 (.LO(net58));
 sky130_fd_sc_hd__conb_1 tiny_user_project_59 (.LO(net59));
 sky130_fd_sc_hd__conb_1 tiny_user_project_60 (.LO(net60));
 sky130_fd_sc_hd__conb_1 tiny_user_project_61 (.LO(net61));
 sky130_fd_sc_hd__conb_1 tiny_user_project_62 (.LO(net62));
 sky130_fd_sc_hd__conb_1 tiny_user_project_63 (.LO(net63));
 sky130_fd_sc_hd__conb_1 tiny_user_project_64 (.LO(net64));
 sky130_fd_sc_hd__conb_1 tiny_user_project_65 (.LO(net65));
 sky130_fd_sc_hd__conb_1 tiny_user_project_66 (.LO(net66));
 sky130_fd_sc_hd__conb_1 tiny_user_project_67 (.LO(net67));
 sky130_fd_sc_hd__conb_1 tiny_user_project_68 (.LO(net68));
 sky130_fd_sc_hd__conb_1 tiny_user_project_69 (.LO(net69));
 sky130_fd_sc_hd__conb_1 tiny_user_project_70 (.LO(net70));
 sky130_fd_sc_hd__conb_1 tiny_user_project_71 (.LO(net71));
 sky130_fd_sc_hd__conb_1 tiny_user_project_72 (.LO(net72));
 sky130_fd_sc_hd__conb_1 tiny_user_project_73 (.LO(net73));
 sky130_fd_sc_hd__conb_1 tiny_user_project_74 (.LO(net74));
 sky130_fd_sc_hd__conb_1 tiny_user_project_75 (.LO(net75));
 sky130_fd_sc_hd__conb_1 tiny_user_project_76 (.LO(net76));
 sky130_fd_sc_hd__conb_1 tiny_user_project_77 (.LO(net77));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_io_in[0]  (.A(io_in[0]),
    .X(clknet_0_io_in[0]));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__dlymetal6s2s_1 input1 (.A(io_in[1]),
    .X(net1));
 sky130_fd_sc_hd__buf_2 output2 (.A(net2),
    .X(io_out[18]));
 sky130_fd_sc_hd__buf_2 output3 (.A(net3),
    .X(io_out[19]));
 sky130_fd_sc_hd__buf_2 output4 (.A(net4),
    .X(io_out[20]));
 sky130_fd_sc_hd__buf_2 output5 (.A(net5),
    .X(io_out[21]));
 sky130_fd_sc_hd__buf_2 output6 (.A(net6),
    .X(io_out[22]));
 sky130_fd_sc_hd__buf_2 output7 (.A(net7),
    .X(io_out[23]));
 sky130_fd_sc_hd__buf_2 output8 (.A(net8),
    .X(io_out[24]));
 sky130_fd_sc_hd__buf_2 output9 (.A(net9),
    .X(io_out[25]));
 sky130_fd_sc_hd__conb_1 tiny_user_project_10 (.LO(net10));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_0__f_io_in[0]  (.A(clknet_0_io_in[0]),
    .X(clknet_2_0__leaf_io_in[0]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_1__f_io_in[0]  (.A(clknet_0_io_in[0]),
    .X(clknet_2_1__leaf_io_in[0]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_2__f_io_in[0]  (.A(clknet_0_io_in[0]),
    .X(clknet_2_2__leaf_io_in[0]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_3__f_io_in[0]  (.A(clknet_0_io_in[0]),
    .X(clknet_2_3__leaf_io_in[0]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\mod._d_io_out[7] ),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\mod._d_io_out[3] ),
    .X(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__186__D (.DIODE(_000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__142__B1 (.DIODE(_000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__133__B1 (.DIODE(_000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__119__B1 (.DIODE(_000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__108__B1 (.DIODE(_000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__159__A2 (.DIODE(_048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__155__C (.DIODE(_048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__184__B1 (.DIODE(_069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__179__A (.DIODE(_069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__176__A (.DIODE(_069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__167__A (.DIODE(_069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__158__A (.DIODE(_069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__103__A (.DIODE(_069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__097__A (.DIODE(_069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__095__B (.DIODE(_069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__094__A (.DIODE(_069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__174__A (.DIODE(_071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__164__A (.DIODE(_071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__155__A (.DIODE(_071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__151__B1 (.DIODE(_071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__131__A (.DIODE(_071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__126__B1 (.DIODE(_071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__125__A (.DIODE(_071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__121__B1 (.DIODE(_071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__102__A (.DIODE(_071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__098__B1 (.DIODE(_071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__181__B1 (.DIODE(_075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__169__B1 (.DIODE(_075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__160__B1 (.DIODE(_075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__149__A (.DIODE(_075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__145__A (.DIODE(_075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__139__A (.DIODE(_075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__136__A (.DIODE(_075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__114__A (.DIODE(_075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__111__A (.DIODE(_075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__105__A (.DIODE(_075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__117__C (.DIODE(_076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__110__C (.DIODE(_076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__108__A2 (.DIODE(_076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__107__B (.DIODE(_076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__105__B (.DIODE(_076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__130__C (.DIODE(_086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__124__C (.DIODE(_086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__123__A2 (.DIODE(_086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__122__A2 (.DIODE(_086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__121__A2 (.DIODE(_086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__120__A (.DIODE(_086_));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_0_io_in[0]_A  (.DIODE(io_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(io_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__195__D (.DIODE(\mod._d_io_out[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__184__A2 (.DIODE(\mod._d_io_out[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__183__A1 (.DIODE(\mod._d_io_out[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__182__A1 (.DIODE(\mod._d_io_out[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__181__A1 (.DIODE(\mod._d_io_out[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__117__B (.DIODE(\mod._q_cnt[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__110__B (.DIODE(\mod._q_cnt[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__108__A1 (.DIODE(\mod._q_cnt[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__107__A (.DIODE(\mod._q_cnt[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__116__B (.DIODE(\mod._q_cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__115__A1 (.DIODE(\mod._q_cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__113__A (.DIODE(\mod._q_cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__093__A (.DIODE(net1));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_297 ();
 assign io_oeb[0] = net41;
 assign io_oeb[10] = net51;
 assign io_oeb[11] = net52;
 assign io_oeb[12] = net53;
 assign io_oeb[13] = net54;
 assign io_oeb[14] = net55;
 assign io_oeb[15] = net56;
 assign io_oeb[16] = net57;
 assign io_oeb[17] = net58;
 assign io_oeb[18] = net59;
 assign io_oeb[19] = net60;
 assign io_oeb[1] = net42;
 assign io_oeb[20] = net61;
 assign io_oeb[21] = net62;
 assign io_oeb[22] = net63;
 assign io_oeb[23] = net64;
 assign io_oeb[24] = net65;
 assign io_oeb[25] = net66;
 assign io_oeb[26] = net67;
 assign io_oeb[27] = net68;
 assign io_oeb[28] = net69;
 assign io_oeb[29] = net70;
 assign io_oeb[2] = net43;
 assign io_oeb[30] = net71;
 assign io_oeb[31] = net72;
 assign io_oeb[32] = net73;
 assign io_oeb[33] = net74;
 assign io_oeb[34] = net75;
 assign io_oeb[35] = net76;
 assign io_oeb[36] = net77;
 assign io_oeb[37] = net10;
 assign io_oeb[3] = net44;
 assign io_oeb[4] = net45;
 assign io_oeb[5] = net46;
 assign io_oeb[6] = net47;
 assign io_oeb[7] = net48;
 assign io_oeb[8] = net49;
 assign io_oeb[9] = net50;
 assign io_out[0] = net11;
 assign io_out[10] = net21;
 assign io_out[11] = net22;
 assign io_out[12] = net23;
 assign io_out[13] = net24;
 assign io_out[14] = net25;
 assign io_out[15] = net26;
 assign io_out[16] = net27;
 assign io_out[17] = net28;
 assign io_out[1] = net12;
 assign io_out[26] = net29;
 assign io_out[27] = net30;
 assign io_out[28] = net31;
 assign io_out[29] = net32;
 assign io_out[2] = net13;
 assign io_out[30] = net33;
 assign io_out[31] = net34;
 assign io_out[32] = net35;
 assign io_out[33] = net36;
 assign io_out[34] = net37;
 assign io_out[35] = net38;
 assign io_out[36] = net39;
 assign io_out[37] = net40;
 assign io_out[3] = net14;
 assign io_out[4] = net15;
 assign io_out[5] = net16;
 assign io_out[6] = net17;
 assign io_out[7] = net18;
 assign io_out[8] = net19;
 assign io_out[9] = net20;
endmodule

